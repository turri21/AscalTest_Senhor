---------------------------------------------------------------------------------
-- ASCAL_TEST
---------------------------------------------------------------------------------

-- A IAUTO
-- B HIMIN
-- C HIMAX
-- D VIMIN
-- E VIMAX
-- F OAUTO
-- G OHMIN
-- H OHMAX
-- I OVMIN
-- J OVMAX
-- K Mire
-- L RESET
-- M Double resolutiuon
-- N Interleaved

-- +/-, O/P
-- ++ / -- , 9/0

--  A,B : IHMIN
--  IHMAX

LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
USE IEEE.numeric_std.all;
USE IEEE.std_logic_unsigned.ALL;

LIBRARY work;
USE work.base_pack.ALL;

ENTITY emu IS
  PORT (
    -- Master input clock
    clk_50m          : IN    std_logic;

    -- Async reset from top-level module. Can be used as initial reset.
    reset            : IN    std_logic;

    -- Must be passed to hps_io module
    hps_bus          : INOUT std_logic_vector(45 DOWNTO 0);

    -- Base video clock. Usually equals to CLK_SYS.
    clk_video        : OUT   std_logic;

    -- Multiple resolutions are supported using different CE_PIXEL rates.
    -- Must be based on CLK_VIDEO
    ce_pixel         : OUT   std_logic;

    -- VGA
    vga_r            : OUT   std_logic_vector(7 DOWNTO 0);
    vga_g            : OUT   std_logic_vector(7 DOWNTO 0);
    vga_b            : OUT   std_logic_vector(7 DOWNTO 0);
    vga_hs           : OUT   std_logic; -- positive pulse!
    vga_vs           : OUT   std_logic; -- positive pulse!
    vga_f1           : OUT   std_logic;
    vga_de           : OUT   std_logic; -- = not (VBlank or HBlank)
    vga_sl           : OUT   std_logic_vector(1 DOWNTO 0);

    -- LED
    led_user         : OUT   std_logic; -- 1 - ON, 0 - OFF.

    -- b[1]: 0 - LED status is system status ORed with b[0]
    --       1 - LED status is controled solely by b[0]
    -- hint: supply 2'b00 to let the system control the LED.
    led_power        : OUT   std_logic_vector(1 DOWNTO 0);
    led_disk         : OUT   std_logic_vector(1 DOWNTO 0);
    
    -- Video aspect ratio for HDMI. Most retro systems have ratio 4:3.
    video_arx        : OUT   std_logic_vector(7 DOWNTO 0);
    video_ary        : OUT   std_logic_vector(7 DOWNTO 0);

    -- AUDIO
    audio_l          : OUT   std_logic_vector(15 DOWNTO 0);
    audio_r          : OUT   std_logic_vector(15 DOWNTO 0);
    audio_s          : OUT   std_logic; -- 1 = signed audio, 0 = unsigned
    -- 0 - no mix, 1 - 25%, 2 - 50%, 3 - 100% (mono)
    audio_mix        : OUT   std_logic_vector(1 DOWNTO 0);

    adc_bus          : INOUT std_logic_vector(3 DOWNTO 0);
    
    tape_in          : IN    std_logic;

    buttons          : IN    std_logic_vector(1 DOWNTO 0);
    
    -- SD-SPI
    sd_sck           : OUT   std_logic := 'Z';
    sd_mosi          : OUT   std_logic := 'Z';
    sd_miso          : IN    std_logic;
    sd_cs            : OUT   std_logic := 'Z';
    sd_cd            : IN    std_logic;
    
    ----------------------------------------------
    sconf   : OUT   std_logic_vector(4 DOWNTO 0);
    
    iauto   : OUT std_logic; -- 1=Autodetect image size 0=Choose window
    himin   : OUT natural RANGE 0 TO 4095;
    himax   : OUT natural RANGE 0 TO 4095;
    vimin   : OUT natural RANGE 0 TO 4095;
    vimax   : OUT natural RANGE 0 TO 4095;
    
    hdisp   : IN  natural RANGE 0 TO 4095;
    hmin    : OUT natural RANGE 0 TO 4095;
    hmax    : OUT natural RANGE 0 TO 4095;
    vdisp   : IN  natural RANGE 0 TO 4095;
    vmin    : OUT natural RANGE 0 TO 4095;
    vmax    : OUT natural RANGE 0 TO 4095;

    ----------------------------------------------
    -- High latency DDR3 RAM interface
    -- Use for non-critical time purposes
    ddram_clk        : OUT   std_logic;
    ddram_busy       : IN    std_logic;
    ddram_burstcnt   : OUT   std_logic_vector(7 DOWNTO 0);
    ddram_addr       : OUT   std_logic_vector(28 DOWNTO 0);
    ddram_dout       : IN    std_logic_vector(63 DOWNTO 0);
    ddram_dout_ready : IN    std_logic;
    ddram_rd         : OUT   std_logic;
    ddram_din        : OUT   std_logic_vector(63 DOWNTO 0);
    ddram_be         : OUT   std_logic_vector(7 DOWNTO 0);
    ddram_we         : OUT   std_logic;

    -- SDRAM interface with lower latency
    sdram_clk        : OUT   std_logic;
    sdram_cke        : OUT   std_logic;
    sdram_a          : OUT   std_logic_vector(12 DOWNTO 0);
    sdram_ba         : OUT   std_logic_vector(1 DOWNTO 0);
    sdram_dq         : INOUT std_logic_vector(15 DOWNTO 0);
    sdram_dqml       : OUT   std_logic;
    sdram_dqmh       : OUT   std_logic;
    sdram_ncs        : OUT   std_logic;
    sdram_ncas       : OUT   std_logic;
    sdram_nras       : OUT   std_logic;
    sdram_nwe        : OUT   std_logic;
    
    uart_cts         : IN    std_logic;
    uart_rts         : OUT   std_logic;
    uart_rxd         : IN    std_logic;
    uart_txd         : OUT   std_logic;
    uart_dtr         : OUT   std_logic;
    uart_dsr         : IN    std_logic;
    
    user_in          : IN    std_logic_vector(5 DOWNTO 0);
    user_out         : OUT   std_logic_vector(5 DOWNTO 0);
    
    osd_status       : IN    std_logic);
END emu;

ARCHITECTURE struct OF emu IS

  COMPONENT pll IS
    PORT (
      refclk   : in  std_logic; -- clk
      rst      : in  std_logic; -- reset
      outclk_0 : out std_logic; -- clk
      outclk_1 : out std_logic; -- clk
      locked   : out std_logic  -- export
      );
  END COMPONENT pll;
  
  CONSTANT CONF_STR : string := 
    "SCALERTEST;;" &
    "O46,Scaler,Nearest,Bilinear,SharpBilinear,Bicubic,Poly,Poly,Poly,TEST;" &
    "O7,Scaler,Direct,TripleBuffer;" &
    "O8,Scaler,Normal,Synchro;" &
    "V1.0";

  FUNCTION to_slv(s: string) return std_logic_vector is 
    CONSTANT ss : string(1 to s'length) := s; 
    VARIABLE rval : std_logic_vector(1 to 8 * s'length); 
    VARIABLE p : integer; 
    VARIABLE c : integer; 
  BEGIN
    FOR i in ss'range LOOP
      p := 8 * i;
      c := character'pos(ss(i));
      rval(p - 7 to p) := std_logic_vector(to_unsigned(c,8)); 
    END LOOP;
    RETURN rval;
  END FUNCTION; 

  COMPONENT hps_io
    GENERIC (
      STRLEN : integer;
      PS2DIV : integer := 1000;
      WIDE   : integer := 0; --  8bits download bus
      VDNUM  : integer := 1;
      PS2WE  : integer := 0);
    PORT (
      clk_sys           : IN  std_logic;
      hps_bus           : INOUT std_logic_vector(45 DOWNTO 0);

      conf_str          : IN  std_logic_vector(8*STRLEN-1 DOWNTO 0);
      joystick_0        : OUT std_logic_vector(31 DOWNTO 0);
      joystick_1        : OUT std_logic_vector(31 DOWNTO 0);
      joystick_2        : OUT std_logic_vector(31 DOWNTO 0);
      joystick_3        : OUT std_logic_vector(31 DOWNTO 0);
      joystick_4        : OUT std_logic_vector(31 DOWNTO 0);
      joystick_5        : OUT std_logic_vector(31 DOWNTO 0);
      joystick_analog_0 : OUT std_logic_vector(15 DOWNTO 0);
      joystick_analog_1 : OUT std_logic_vector(15 DOWNTO 0);
      joystick_analog_2 : OUT std_logic_vector(15 DOWNTO 0);
      joystick_analog_3 : OUT std_logic_vector(15 DOWNTO 0);
      joystick_analog_4 : OUT std_logic_vector(15 DOWNTO 0);
      joystick_analog_5 : OUT std_logic_vector(15 DOWNTO 0);
      buttons           : OUT std_logic_vector(1 DOWNTO 0);
      forced_scandoubler: OUT std_logic;
      status            : OUT std_logic_vector(31 DOWNTO 0);
      status_in         : IN  std_logic_vector(31 DOWNTO 0);
      status_set        : IN  std_logic;
      status_menumask   : IN  std_logic_vector(15 DOWNTO 0);
      new_vmode         : IN  std_logic;
      img_mounted       : OUT std_logic;
      img_readonly      : OUT std_logic;
      img_size          : OUT std_logic_vector(63 DOWNTO 0);
      sd_lba            : IN  std_logic_vector(31 DOWNTO 0);
      sd_rd             : IN  std_logic;
      sd_wr             : IN  std_logic;
      sd_ack            : OUT std_logic;
      sd_conf           : IN  std_logic;
      sd_ack_conf       : OUT std_logic;
      sd_buff_addr      : OUT std_logic_vector(8 DOWNTO 0);
      sd_buff_dout      : OUT std_logic_vector(7 DOWNTO 0);
      sd_buff_din       : IN  std_logic_vector(7 DOWNTO 0);
      sd_buff_wr        : OUT std_logic;
      ioctl_download    : OUT std_logic;
      ioctl_index       : OUT std_logic_vector(7 DOWNTO 0);
      ioctl_wr          : OUT std_logic;
      ioctl_addr        : OUT std_logic_vector(24 DOWNTO 0);
      ioctl_dout        : OUT std_logic_vector(7 DOWNTO 0);
      ioctl_wait        : IN  std_logic;
      rtc               : OUT std_logic_vector(64 DOWNTO 0);
      timestamp         : OUT std_logic_vector(32 DOWNTO 0);
      uart_mode         : IN  std_logic_vector(15 DOWNTO 0);
      ps2_kbd_clk_out   : OUT std_logic;
      ps2_kbd_data_out  : OUT std_logic;
      ps2_kbd_clk_in    : IN  std_logic;
      ps2_kbd_data_in   : IN  std_logic;
      ps2_kbd_led_use   : IN  std_logic_vector(2 DOWNTO 0);
      ps2_kbd_led_status: IN  std_logic_vector(2 DOWNTO 0);
      ps2_mouse_clk_out : OUT std_logic;
      ps2_mouse_data_out: OUT std_logic;
      ps2_mouse_clk_in  : IN  std_logic;
      ps2_mouse_data_in : IN  std_logic;
      ps2_key           : OUT std_logic_vector(10 DOWNTO 0);
      ps2_mouse         : OUT std_logic_vector(24 DOWNTO 0);
      ps2_mouse_ext     : OUT std_logic_vector(15 DOWNTO 0));
  END COMPONENT hps_io;

  SIGNAL status          : std_logic_vector(31 DOWNTO 0);
  SIGNAL status_in       : std_logic_vector(31 DOWNTO 0):=x"00000000";
  SIGNAL status_set      : std_logic :='0';
  SIGNAL status_menumask : std_logic_vector(15 DOWNTO 0):=x"0000";
  SIGNAL new_vmode       : std_logic :='0';

  SIGNAL ioctl_wait : std_logic :='0';
  
  SIGNAL ps2_key,ps2_key_delay : std_logic_vector(10 DOWNTO 0);
  SIGNAL key_0,key_1,key_2,key_3,key_4,key_5,key_6,key_7,key_8,key_9 : std_logic;
  SIGNAL key_a,key_b,key_c,key_d,key_e,key_f,key_g,key_h,key_i,key_j : std_logic;
  SIGNAL key_k,key_l,key_m,key_n,key_o,key_p,key_q,key_r,key_s,key_t : std_logic;
  SIGNAL key_u,key_v,key_w,key_x,key_y,key_z                         : std_logic;
  SIGNAL key_space,key_return                                        : std_logic;
  
  SIGNAL clksys,clksys2,pll_locked : std_logic;
  
  SIGNAL reset_na : std_logic;
  
  ------------------------------------------------
  SIGNAL sel : natural RANGE 0 TO 10;
  SIGNAL mire : natural RANGE 0 TO 15 := 0;
  SIGNAL iauto_n_i : std_logic :='0';
  SIGNAL oauto_n_i : std_logic :='0';
  SIGNAL inc,dec : std_logic;
  SIGNAL delta : natural RANGE 1 TO 10;
  SIGNAL double : std_logic :='0';
  
  ------------------------------------------------
  SIGNAL gde,ghs,gvs,gce : std_logic;
  SIGNAL gfl : std_logic :='0';
  SIGNAL inter : std_logic :='0';
  SIGNAL ghcpt,gvcpt : natural RANGE 0 TO 4095;
  CONSTANT CGHDISP : natural :=640; --320; --120; --1440; --374; --320; --640; --160;
  CONSTANT CGVDISP : natural :=400; --287; --256; --256; --400; --100;
  
  SIGNAL ghdisp      : natural range 0 to 4095 := CGHDISP; --640; --320; --800;
  SIGNAL ghsyncstart : natural range 0 to 4095 := CGHDISP+88;
  SIGNAL ghsyncend   : natural range 0 to 4095 := CGHDISP+88+48;
  SIGNAL ghtotal     : natural range 0 to 4095 := CGHDISP+88+48+40;
  
  SIGNAL gvdisp      : natural range 0 to 4095 := CGVDISP; --400; --600;
  SIGNAL gvsyncstart : natural range 0 to 4095 := CGVDISP+1;
  SIGNAL gvsyncend   : natural range 0 to 4095 := CGVDISP+1+4;
  SIGNAL gvtotal     : natural range 0 to 4095 := CGVDISP+1+4+20;
  SIGNAL gr,gg,gb    : uv8;
  SIGNAL calt : natural RANGE 0 TO 63;

  SIGNAL move, dir : std_logic;
  SIGNAL clkdiv : uint24;
  ------------------------------------------------
  SIGNAL himin_i : natural RANGE 0 TO 4095 := 0;
  -- 315 313 312  .311.  310 309 308 307
  SIGNAL himax_i : natural RANGE 0 TO 4095 := 319; --306; --251; --CGHDISP-1;
  SIGNAL vimin_i : natural RANGE 0 TO 4095 := 0;
  SIGNAL vimax_i : natural RANGE 0 TO 4095 :=CGVDISP-1;
  SIGNAL hmin_i,hmax_i : natural RANGE 0 TO 4095;
  SIGNAL vmin_i,vmax_i : natural RANGE 0 TO 4095;
  
  -- OVO -----------------------------------------
  FUNCTION CC(i : character) RETURN unsigned IS
  BEGIN
    CASE i IS
      WHEN '0' => RETURN "00000";
      WHEN '1' => RETURN "00001";
      WHEN '2' => RETURN "00010";
      WHEN '3' => RETURN "00011";
      WHEN '4' => RETURN "00100";
      WHEN '5' => RETURN "00101";
      WHEN '6' => RETURN "00110";
      WHEN '7' => RETURN "00111";
      WHEN '8' => RETURN "01000";
      WHEN '9' => RETURN "01001";
      WHEN 'A' => RETURN "01010";
      WHEN 'B' => RETURN "01011";
      WHEN 'C' => RETURN "01100";
      WHEN 'D' => RETURN "01101";
      WHEN 'E' => RETURN "01110";
      WHEN 'F' => RETURN "01111";
      WHEN ' ' => RETURN "10000";
      WHEN '=' => RETURN "10001";
      WHEN '+' => RETURN "10010";
      WHEN '-' => RETURN "10011";
      WHEN '<' => RETURN "10100";
      WHEN '>' => RETURN "10101";
      WHEN '^' => RETURN "10110";
      WHEN 'v' => RETURN "10111";
      WHEN '(' => RETURN "11000";
      WHEN ')' => RETURN "11001";
      WHEN ':' => RETURN "11010";
      WHEN '.' => RETURN "11011";
      WHEN ',' => RETURN "11100";
      WHEN '?' => RETURN "11101";
      WHEN '|' => RETURN "11110";
      WHEN '#' => RETURN "11111";
      WHEN OTHERS => RETURN "10000";
    END CASE;
  END FUNCTION CC;
  FUNCTION CS(s : string) RETURN unsigned IS
    VARIABLE r : unsigned(0 TO s'length*5-1);
    VARIABLE j : natural :=0;
  BEGIN
    FOR i IN s'RANGE LOOP
      r(j TO j+4) :=CC(s(i));
      j:=j+5;
    END LOOP;
    RETURN r;
  END FUNCTION CS;
  FUNCTION CN(v : unsigned) RETURN unsigned IS
    VARIABLE t : unsigned(0 TO v'length-1);
    VARIABLE o : unsigned(0 TO v'length/4*5-1);
  BEGIN
    t:=v;
    FOR i IN 0 TO v'length/4-1 LOOP
      o(i*5 TO i*5+4):='0' & t(i*4 TO i*4+3);
    END LOOP;
    RETURN o;
  END FUNCTION CN;

  ------------------------------------------------
  SIGNAL vga_r_u   : unsigned(7 DOWNTO 0);
  SIGNAL vga_g_u   : unsigned(7 DOWNTO 0);
  SIGNAL vga_b_u   : unsigned(7 DOWNTO 0);
  
  -- OVO -----------------------------------------
  SIGNAL ovo_ena  : std_logic;
  SIGNAL ovo_in0  : unsigned(0 TO 32*5-1) :=(OTHERS =>'0');
  SIGNAL ovo_in1  : unsigned(0 TO 32*5-1) :=(OTHERS =>'0');
  
  ------------------------------------------------
  CONSTANT test : unsigned(0 TO 320*128-1):=
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000111000000000000000000000000000000000011111000011100001110011100111111100011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000001111000001110000111001110011111110001111000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000001000000000000000000000000000000000000100000000100000100001000100100100100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000010000000000000000000000000000010000100000010000010000100010010010010000100000000000000000000000000000000000000000000000000000000000000000000000" &
"00000010100000000000000011000000000000000000100000001010000100001000100100101000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000010000000000000110000000000000100000010000101000010000100010010010100000010000000000000000000000000000000000000000000000000000000000000000000000" &
"00000010100000000000000011000000000000000000100000001010000100001000000100001000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000110000000000000100000010000101000010000100000010000100000010000000000000000000000000000000000000000000000000000000000000000000000" &
"00000100010000000000000000000000000000000000100000010001000100001000000100001000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000100000010001000100010000100000010000100000010000000000000000000000000000000000000000000000000000000000000000000000" &
"00000111110000000000000000000000000000000000100000011111000100001000000100001000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000100000010001111100010000100000010000100000010000000000000000000000000000000000000000000000000000000000000000000000" &
"00001000001000000000000000000000000000000000100000100000100100001000000100001000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000100000010010000010010000100000010000100000010000000000000000000000000000000000000000000000000000000000000000000000" &
"00001000001000000000000011000000000000000000100000100000100100001000000100000100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000110000000000000010000100010000010010000100000010000010000100000000000000000000000000000000000000000000000000000000000000000000000" &
"00011110111100000000000011000000000000000011111001111011110011110000011111000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000110000000000000001111000111101111001111000001111100001111000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00001111110000000000000000000000000000000111010000000000000111000000000000000000000000100000000000000011100111000111110011100011100111110011100111000000000000000000000000001110100000000000000000000000000000001110100000000000001110000000000000000000000001000000000000000001111000111001110111000111001111100111001110000000" &
"00000100001000000000000000000000000000001000110000000000000001000000000000000000000000100000000000000001000010000001000001100011000001000001100010000000000000000000000000010001100000000000000000000000000000010001100000000000000010000000000000000000000001000000000000000010000100010000100011000110000010000011000100000000" &
"00000100001000000000000011000000000000001000010000011100000001000000011100000011101001111100000000000001000010000001000001010111000001000001010010000000000000000000000000100000100000000000000110000000000000010000100000111000000010000000111000000111010011111000000000000100000010010000100010101110000010000010100100000000" &
"00000100001000000000000011000000000000001000000000100010000001000000100010000100011000100000000000000001000010000001000001010101000001000001010010000000000000000000000000100000000000000000000110000000000000010000000001000100000010000001000100001000110001000000000000000100000010010000100010101010000010000010100100000000" &
"00000111110000000000000000000000000000000111100001000001000001000001000001001000001000100000000000000001111110000001000001001001000001000001001010000000000000000000000000100000000000000000000000000000000000001111000010000010000010000010000010010000010001000000000000000100000010011111100010010010000010000010010100000000" &
"00000100001000000000000000000000000000000000010001111111000001000001111111001000000000100000000000000001000010000001000001001001000001000001001010000000000000000000000000100011110000000000000000000000000000000000100011111110000010000011111110010000000001000000000000000100000010010000100010010010000010000010010100000000" &
"00000100001000000000000000000000000000001000010001000000000001000001000000001000000000100000000000000001000010000001000001000001000001000001000110000000000000000000000000100000100000000000000000000000000000010000100010000000000010000010000000010000000001000000000000000100000010010000100010000010000010000010001100000000" &
"00000100001000000000000011000000000000001100010000100001000001000000100001000100001000100010000000000001000010000001000001000001000001000001000110000000000000000000000000010000100000000000000110000000000000011000100001000010000010000001000010001000010001000100000000000010000100010000100010000010000010000010001100000000" &
"00001111110000000000000011000000000000001011100000011110000111110000011110000011110000011100000000000011100111000111110011100011100111110011100010000000000000000000000000001111000000000000000110000000000000010111000000111100001111100000111100000111100000111000000000000001111000111001110111000111001111100111000100000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000011101000000000000000000000000000000111010000000000000111000000000000000000000000100000000000000011100111000111110011100011100111000011100111000000000000000000000000111001110000000000000000000000000000001110100000000000001110000000000000000000000001000000000000000001111000111001110111000111001110000111001110000000" &
"00000100011000000000000000000000000000001000110000000000000001000000000000000000000000100000000000000001000010000001000001100011000001000001000010000000000000000000000000010000100000000000000000000000000000010001100000000000000010000000000000000000000001000000000000000010000100010000100011000110000010000010000100000000" &
"00001000001000000000000011000000000000001000010000011100000001000000011100000011101001111100000000000001000010000001000001010111000010100000100100000000000000000000000000010000100000000000000110000000000000010000100000111000000010000000111000000111010011111000000000000100000010010000100010101110000101000001001000000000" &
"00001000000000000000000011000000000000001000000000100010000001000000100010000100011000100000000000000001000010000001000001010101000010100000100100000000000000000000000000010000100000000000000110000000000000010000000001000100000010000001000100001000110001000000000000000100000010010000100010101010000101000001001000000000" &
"00001000000000000000000000000000000000000111100001000001000001000001000001001000001000100000000000000001111110000001000001001001000100010000011000000000000000000000000000011111100000000000000000000000000000001111000010000010000010000010000010010000010001000000000000000100000010011111100010010010001000100000110000000000" &
"00001000000000000000000000000000000000000000010001111111000001000001111111001000000000100000000000000001000010000001000001001001000111110000100100000000000000000000000000010000100000000000000000000000000000000000100011111110000010000011111110010000000001000000000000000100000010010000100010010010001111100001001000000000" &
"00001000000000000000000000000000000000001000010001000000000001000001000000001000000000100000000000000001000010000001000001000001001000001000100100000000000000000000000000010000100000000000000000000000000000010000100010000000000010000010000000010000000001000000000000000100000010010000100010000010010000010001001000000000" &
"00000100001000000000000011000000000000001100010000100001000001000000100001000100001000100010000000000001000010000001000001000001001000001001000010000000000000000000000000010000100000000000000110000000000000011000100001000010000010000001000010001000010001000100000000000010000100010000100010000010010000010010000100000000" &
"00000011110000000000000011000000000000001011100000011110000111110000011110000011110000011100000000000011100111000111110011100011111110111111100111000000000000000000000000111001110000000000000110000000000000010111000000111100001111100000111100000111100000111000000000000001111000111001110111000111111101111111001110000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00011111100000000000000000000000000000000111010000000000000111000000000000000000000000100000000000000011100011100111110011100011100111110011100111000000000000000000000000001111100000000000000000000000000000001110100000000000001110000000000000000000000001000000000000000001111000111000111111000111001111100111001110000000" &
"00001000010000000000000000000000000000001000110000000000000001000000000000000000000000100000000000000001000001000001000001100011000001000001100010000000000000000000000000000010000000000000000000000000000000010001100000000000000010000000000000000000000001000000000000000010000100010000010011000110000010000011000100000000" &
"00001000001000000000000011000000000000001000010000011100000001000000011100000011101001111100000000000001000001000001000001010111000001000001010010000000000000000000000000000010000000000000000110000000000000010000100000111000000010000000111000000111010011111000000000000100000010010000010010101110000010000010100100000000" &
"00001000001000000000000011000000000000001000000000100010000001000000100010000100011000100000000000000000100010000001000001010101000001000001010010000000000000000000000000000010000000000000000110000000000000010000000001000100000010000001000100001000110001000000000000000100000010001000100010101010000010000010100100000000" &
"00001000001000000000000000000000000000000111100001000001000001000001000001001000001000100000000000000000100010000001000001001001000001000001001010000000000000000000000000000010000000000000000000000000000000001111000010000010000010000010000010010000010001000000000000000100000010001000100010010010000010000010010100000000" &
"00001000001000000000000000000000000000000000010001111111000001000001111111001000000000100000000000000000010100000001000001001001000001000001001010000000000000000000000000000010000000000000000000000000000000000000100011111110000010000011111110010000000001000000000000000100000010000101000010010010000010000010010100000000" &
"00001000001000000000000000000000000000001000010001000000000001000001000000001000000000100000000000000000010100000001000001000001000001000001000110000000000000000000000000000010000000000000000000000000000000010000100010000000000010000010000000010000000001000000000000000100000010000101000010000010000010000010001100000000" &
"00001000010000000000000011000000000000001100010000100001000001000000100001000100001000100010000000000000001000000001000001000001000001000001000110000000000000000000000000000010000000000000000110000000000000011000100001000010000010000001000010001000010001000100000000000010000100000010000010000010000010000010001100000000" &
"00011111100000000000000011000000000000001011100000011110000111110000011110000011110000011100000000000000001000000111110011100011100111110011100010000000000000000000000000001111100000000000000110000000000000010111000000111100001111100000111100000111100000111000000000000001111000000010000111000111001111100111000100000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00001111111000000000000000000000000000000111010000000000000111000000000000000000000000100000000000000011100011100111110011100011100111000011100111000000000000000000000000000111110000000000000000000000000000001110100000000000001110000000000000000000000001000000000000000001111000111000111111000111001110000111001110000000" &
"00000100001000000000000000000000000000001000110000000000000001000000000000000000000000100000000000000001000001000001000001100011000001000001000010000000000000000000000000000001000000000000000000000000000000010001100000000000000010000000000000000000000001000000000000000010000100010000010011000110000010000010000100000000" &
"00000100001000000000000011000000000000001000010000011100000001000000011100000011101001111100000000000001000001000001000001010111000010100000100100000000000000000000000000000001000000000000000110000000000000010000100000111000000010000000111000000111010011111000000000000100000010010000010010101110000101000001001000000000" &
"00000100100000000000000011000000000000001000000000100010000001000000100010000100011000100000000000000000100010000001000001010101000010100000100100000000000000000000000000000001000000000000000110000000000000010000000001000100000010000001000100001000110001000000000000000100000010001000100010101010000101000001001000000000" &
"00000111100000000000000000000000000000000111100001000001000001000001000001001000001000100000000000000000100010000001000001001001000100010000011000000000000000000000000000000001000000000000000000000000000000001111000010000010000010000010000010010000010001000000000000000100000010001000100010010010001000100000110000000000" &
"00000100100000000000000000000000000000000000010001111111000001000001111111001000000000100000000000000000010100000001000001001001000111110000100100000000000000000000000000010001000000000000000000000000000000000000100011111110000010000011111110010000000001000000000000000100000010000101000010010010001111100001001000000000" &
"00000100001000000000000000000000000000001000010001000000000001000001000000001000000000100000000000000000010100000001000001000001001000001000100100000000000000000000000000010001000000000000000000000000000000010000100010000000000010000010000000010000000001000000000000000100000010000101000010000010010000010001001000000000" &
"00000100001000000000000011000000000000001100010000100001000001000000100001000100001000100010000000000000001000000001000001000001001000001001000010000000000000000000000000010001000000000000000110000000000000011000100001000010000010000001000010001000010001000100000000000010000100000010000010000010010000010010000100000000" &
"00001111111000000000000011000000000000001011100000011110000111110000011110000011110000011100000000000000001000000111110011100011111110111111100111000000000000000000000000001110000000000000000110000000000000010111000000111100001111100000111100000111100000111000000000000001111000000010000111000111111101111111001110000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000011110000000000000001111100000000000000000011110001100001000111100000000000001111100001111110000111100000000000000000000000000000000000000000000000000000000000000000001111000000000000000011110000000000000000001111000110000100011110000000000000111110000111111000011110000000000011000000111000000000000000000000000000" &
"00000100001000000000000001000010000000000000000001000001010001001000000000000000001000010001000000001000000000000000000000000000000000000000000000000000000000000000000000010000100000000000000100001000000000000000000100000101000100100000000000000000100001000100000000100000000000000101000001000100000000000000000000000000" &
"00000100001000000000100001000010000000110000000001000001001001010000000000000000001000001001000000010000000000000000000000000000000000000000000000000000000000000000000000010000100000000010000100001000000011000000000100000100100101000000000000000000100000100100000001000000000000001001000010000010000000000000000000000000" &
"00000100001000000001000001000010000000110000000001000001000101010000000000000100001000001001000000010000000000000000000000000000000000000000000000000000000000000000000000010000100000000100000100011000000011000000000100000100010101000000000000010000100000100100000001000000000000000001000010000010000000000000000000000000" &
"00000100001000000010000001111100000000000000000001000001000011010000000000001000001000001001111000010000000000000000000000000000000000000000000000000000000000000000000000001111100000001000000101101000000000000000000100000100001101000000000000100000100000100111100001000000000000000001000010000010000000000000000000000000" &
"00000100001000000100000001000000000000000000000001000001000001010000000000010000001000001001000000010000000000000000000000000000000000000000000000000000000000000000000000000000100000010000000110001000000000000000000100000100000101000000000001000000100000100100000001000000000000000001000010000010000000000000000000000000" &
"00000100001000001000000001000000000000110000000001000001000001010000000000100000001000001001000000010000000000000000000000000000000000000000000000000000000000000000000000000001000000100000000100001000000011000000000100000100000101000000000010000000100000100100000001000000000000000001000010000010000000000000000000000000" &
"00000100001000000000000001000000000000110000000001000001000001001000000000000000001000010001000000001000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000100001000000011000000000100000100000100100000000000000000100001000100000000100000000000000001000001000100000000000000000000000000" &
"00000011110000000000000001000000000000000000000011100001000001000111100000000000001111100001111110000111100000000000000000000000000000000000000000000000000000000000000000001100000000000000000011110000000000000000001110000100000100011110000000000000111110000111111000011110000000000111110000111000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00011101110000000000000000000000000000000011101001000000000000000000000000000000000000000000000000000000000000000000000000100000000100000000000000000000000000000000000000111110000000000000000000000000000000111111000011111110001110100011111110011111110000000000000000000000000000000000000000000000000000000000000000000000" &
"00001000100000000000000000000000000000000100011001000000000000000000000000000000000000000000000000000000000000000000000000100000000100000000000000000000000000000000000000001000000000000000000000000000000000010000100001000010010001100001000010010010010000000000000000000000000000000000000000000000000000000000000000000000" &
"00001001000000000000000011000000000000001000001001011100000111100011011100000111011000011100000000000011011100000111100001111100001111100000011100001100110011011100000000001000000000000000000110000000000000010000100001000010010000100001000010010010010000000000000000000000000000000000000000000000000000000000000000000000" &
"00001010000000000000000011000000000000001000000001100010001000010001100010001000110000100010000000000001100010001000010000100000000100000000100010000101001001100010000000001000000000000000000110000000000000010000100001001000010000000001001000000010000000000000000000000000000000000000000000000000000000000000000000000000" &
"00001110000000000000000000000000000000001000000001000010000000010001000010010000010001000001000000000001000001000000010000100000000100000001000001000110000001000010000000001000000000000000000000000000000000010001000001111000001111000001111000000010000000000000000000000000000000000000000000000000000000000000000000000000" &
"00001001000000000000000000000000000000001000000001000010000111110001000010010000010001111111000000000001000001000111110000100000000100000001111111000100000001000010000000001000010000000000000000000000000000011110000001001000000000100001001000000010000000000000000000000000000000000000000000000000000000000000000000000000" &
"00001000100000000000000000000000000000001000000001000010001000010001000010010000010001000000000000000001000001001000010000100000000100000001000000000100000001000010000000001000010000000000000000000000000000010001000001000010010000100001000010000010000000000000000000000000000000000000000000000000000000000000000000000000" &
"00001000100000000000000011000000000000000100001001000010001000110001000010001000110000100001000000000001100010001000110000100010000100010000100001000100000001000010000000001000010000000000000110000000000000010000100001000010011000100001000010000010000000000000000000000000000000000000000000000000000000000000000000000000" &
"00011100011000000000000011000000000000000011110011100111000111011011100111000111010000011110000000000001011100000111011000011100000011100000011110001111000011100111000000111111110000000000000110000000000000111000010011111110010111000011111110001111100000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000100000000000011110000000000000000001110100000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000100000001000100001000000000000000010001100000000000000000000000001000000000000000000000000000100000100000000000111111100000000000000000000000000000000000000100000100000000011100010000100111111100011111110011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000100000010000000001000001100000000100000100000111100001101110000011111000000000000000000000000110001100000000000000000100000000000000000000000000000000000000110000100000000001000011000100000100000010000000010000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000100000100000000001000001100000000100000000001000010000110001000001000000000000000000000000000101010100001100000000001000001111000011110000111111000000000000101100100011000001000010100100000100000010000000010000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000100001000000000010000000000000000100000000001000010000100001000001000000000000000000000000000100100100001100000000010000010000100100001001001001000000000000100110100011000001000010010100000100000011110000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000100010000000000100000001100000000100000000001000010000100001000001000000000000000000000000000100000100000000000000100000010000100100001001001001000000000000100001100000000001000010001100000100000010000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000100100000000001000000001100000000100000000001000010000100001000001000000000000000000000000000100000100001100000001000000010000100100001001001001000000000000100000100011000001000010000100000100000010000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000100000000000111111000000000000000010000100001000010000100001000001000100000000000000000000000100000100001100000010000000010000100100001001001001000000000000100000100011000001000010000100000100000010000000010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000001111000000111000001110011100000111000000000000000000000000100000100000000000111111000001111000011110001001001000000000000100000100000000011100010000100000100000011111110010000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

  CONSTANT dragon : unsigned(0 TO 260*400-1):= 
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011101110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001101010011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110101101100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000010110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110011011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001101101100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110101110111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111010010111110111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010010111011011010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011101011011111011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110101001111011111011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011010101111011011010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110100110101101101101101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011010011011110111110110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110101110110111110111101101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011101010011111110110101010110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110101111111110111011110111010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011101011010110111101110111010110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111001101111011110110110101011010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001011111011111011011010110110010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001101101111011111110111011011010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101111111110110110011010110010110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000100111011011011111011110110011011010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000001000101111111110110110110111010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000010010111110110111011111010101010110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000010010111011111110110110110110110010110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000100100111111011011110110110101011010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000001001011011010111110101101010110100110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000010101010111111101101110110110100110010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000010010111011011110110101101010110101101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000100101101101101011101101101101010100100101000000000000000000000000000000000000000000000000000000000000000000000000000000010111111110100000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000001000101010111111101111010101010100101101010000000000000000000000000000000000000000000000000000000000000000000000000011111110100000000000100000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000001001011111011011011010101101101010100101001000000000000000000000000000000000000000000000000000000000000000000101111110010000000000001010000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000010010101010110110110111011010101001010100101000000000000000000000000000000000000000000000000000000000010101111110010000000101101111110100000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000100101110101011110110101010011001010101001001000000000000000000000000000000000000000000000000000010111111110100001000110111010110101011100000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000001010101011011110110110110111010101010010101000000000000000000000000000000000000000000000000001011111110100000001000111011011111011101110000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000001000110101101011010101010100101010101001001010100000000000000000000000000000000000000000011111110100000000101010111011110110101101111100000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000010001010110110101101101101010010100100100100010000000000000000000000000000000000000001111110110001000101011010111101101101111111110111000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000100101101111011111011101101101100110010010010100100000000000000000000000000000000011111010100000100110101101111101011111111110101011110000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000101010110101010011011010101010010000100100100000000000000000000000000000000001111111101000001010101011011011101111110110110111111111101000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000001000101011011011011110110101001001101001000100101000000000000000000000000101111101000000010101011011110111111011011011111111101111101100000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000010010101101101101010100101010010100001010001001000010000000000000000000111111100000001010101111101111011110111111101110110101111010111000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000010001011010101011101101100101010010101000000000000000000000000000001111110100000101101011011010111101111111110110111011111111011111111000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000100101010110110100111011010101010010010010000100000000000000000001111110010000010100101101111011110111101101111111101111011011110111010000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000001000110111010101010101010011001001000100000100000000000000000011111110001000010110111110111101111111111011111101101111101110111011101110000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000001010101001101010101010110100101001001000000000000000000000011111101000010011011011011011110111111011101111110111111011011111111111111100000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000010010101101010101010101100110010001000001001000000000000011111010000001011011111101111111111110110111111110111111011111111011101011101000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000101010101010101010101011001001000100000010000000000000101111010000101011011101101111101101111011111110110111111101110110111110111110111000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000100010101010101010010010101010100100100000000000000011111101000010010101101111111101111111101111011011111110110111111101101011101111110000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000001010110101010100100000000010000000000000000000000001111011010001011101111111101101111110110111101111111011011111111010111111111110110100000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000010100101010000000101011011001001000010000000000001111110100000011010111010101111111110111111111111101101101111101101111110110110111111100000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000001001001000111111101101011011001011000000000000111111010000111011111101111111101110111111011110110110111111101111111111011111111101101100000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000110000101111101101001011001011011010010110010000111010000010011111011111101110111011110111110111110111101010111010110101111101101110111000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000100011111101101101101101011001001010010010100100000010101011111011111011111111111111111101011110011010110111011111111111101111111011111000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000011111110110110100100101001011011010110100100100100100010111101111101111101101101110110111110111011011010101101101011101111110111111010000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000011110110010010010100101001001011001010100101101101001000000011111111111101110111111011011011011011010101011011011101110111011011101101110000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000001111011011011010010010100100101001010010110101001001001001000100111101011111111110110111111101101101001000101001101101111111111110111111010000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000111011011001001010010000100001001011001010110111011101011010011000001011111011010111101110110110111010000010000101010110110101101111110101110000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000011101101101001010000000100000100000000011010110101101011011010010001000011011101111101111110110101010101011111100001010011011011110101011111100000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000001111110110000101000010110111101000000000000010101111011111110110110110011000111111101101010110110111010001110101111000001010111110111111111010100000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000111110110010100000001010101000100000000000001111000000111101010110100110100001001011101101101010101001001001111011111111110011010110110101011101100000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000001111011010010000101101010100110100100000001111110010010000111111110111101100110000101101101101110100101000011111100101100111101011101111011101110100000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000111101001000000011010101101010101000000000111111000010101010001111101101101001100010001101101010100110000001111011101111111111101101110101101110111000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000001110100100000010101110110101010000100000001111010010101110111010001111111011111001100010011010101010000010111101100011101101111101010111011011101010100000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000111110110100101010110011010101010101000000111101001001101111010101000011111011010011000100000101001000011111110110011111010111010001101010101101111011000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000001111010010000100011011010101001010000000000111110000101111011111111101000111111011011001000010010000011111110111011111110110100100001011011011101010101000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000111101001000001000101001101010101000000000011110000110111011110110101101101001011110100101001000000111111111011110111101010100100000101101011101101110111000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000001101100100000000101010110101010000101000000010010100101101110111111111011011000111010111111010000101111111011110111110111010000000101001010110101010110101000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000011010010000000001001011010101001010000000001111010001111011101111011101111110110000111111111111111011011110111111101010100000001010000001101011010110011010000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000111101000000000010010101010101100000100000001000000111011110111101111111111011010101111111010101011110111011110110110101000001010000011001010101011010110101000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000001110100000000000101001011010100101010000000011100011001101011110111011011101111110001111110110011101000000111101101011000010010100000101001010110100101011011000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000011110000000000001100101010101010010000000000110000101010010101011110111101111101001011111011001111010000100001011011100110001101000111110010101010101101010101000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000111001000000000001100101010101010100000000001101001010000000001010101110111011101100111111100101110100011111101110110111000011010011111100010100101010101010010000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000001110100000000000011010101010101010000100000011010001110111111101001111101101010101010111110101011111001110000100010101000000110000111101000010010101010101011011000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000011110000000000000111001010101010001010000000101000101010000111110100010110110110110100111101010111100101000000110100010010001101011100011110101010100010100101001000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000111000000000000000110101101101010100100000001110000101011000001011110011011010100100011111011001111010001111000011110110000011010011010001110010010101010101101010000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000001110100000000000001111010101010101010000000000101001010111110000111011100110101000100111110110110111010101111100010111101000111000110110000110001010100101001010011000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000011010000000000000011100101010101000000000000011000001010111110001000111010010100100011111111011011111100001100000011110000000110100100111000011000101001010101010101000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000101100000000000000011011110111000101001000000110100010100101111100011101110101010011011111010100111110011000100000011000101001100001000111000010101000010010010100101000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000110000000000000000111010101001010100010000000101000101010111011100000011011001000011001011111011011101100001110000011010000011010011100011000011000110101001010010100000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000100000000000000001110101101010101001000000011010001010010101111010000110111110010000100101010101111010010000111110110001000010100010100001100100001000010100100100101100000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000001100111101001010000000000010100000101000111011110001001111111001000110010101110101101100100111111100100001101000111110001100000100010100001000010000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000011101010110100001010000000101000101001010101101011000011001111111100011001010011111101001000111111000010010010001100110000100010010000000100101001011000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000110101111100101010000010000110000100101010111011101000010011011111100001100101101100110100001111100101000010000011001011000100000000101001010000100000100000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000111010101010100001010000001100010101010100101010011100100111111011110010110010110011001001000100010000001010001111001011010000101001000000000101001010000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000001110101110101001100000000010010001010101010101101010010000100110111110001100011000100010100000001001000010000011110101100011010111101000100100000000100100000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000011001011101101010001010000011000101010101000101001000100000100110110110000011000110001000010001100100001010001111001100101000010000111111010001001001000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000011101110111100000010000000100000101010100110101010001000001001100110111000111000101100010000010010000010000011111000110100010000110000001111100000000000100000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000110101011101011010000000001010001001010100000010000110110000001100110111000011100010001001000100100001001001111101000010110101110101000000000111110100000001000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000001110111110111100100100000001100100101001010010001111111111000001001101111001011100011100000000010000001000011111011000001110011110110011100000000011101010000000000000000001010000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000001101010111101010010000010011000011010101001000111111111101000010001101111100000110000111100010001001000000111100011001000101010010101001011101001000011101000000000000000010000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000011101011101010101000000000010100100100100100001111111010010000000001001010000011111000001011000100000110001111000000000001110000000011001111011110100000111101000000000001110000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000011010110111111010100001000101000101010010010110110100000000000000010001111100000011100000000010000010000011110100000000001110000000011101011101011011010000011000000001011000000000001010000000000000000000000000000000000" &
"00000000000000000000000000000000000000000111011111111010101000000001010001010101000001010010000101101110000100011111100001111110000001001000001000011101100000100001100000100111000000000101101101001000100010101100000000001010000000000000000000000000000000000000" &
"00000000000000000000000000000000000000001110101011010111000100100001100000101000101011000000101010110111000000111101000000001111101010000001000001111000010100000000000100000110100000000000000010110100010010110000000001011000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000001110111111111010101000000010000101010100000101010101011011111011000001111111110001110101111111010000010001111000100000000000000000000111000000000000000000001011011111101011101111000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000011101010101010110000000100101100010001001011010000101111101101111110011110101010000000110110100000010000001110000000010101010000000001110100011101000000000000000101010111101111000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000011010101111111010101000000010000101010000110100000111110111111101110111011111110000011001100000100000100011110000001000000000000010000101000110110110100010101101010111010110000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000110101011101010101000001000110000100100011001000010111011110110111101111111111111000000010000100000000000111100000100000000000001000001011000101111111111000000010101000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000001111001110111101010100000001010010010001010100001010111111111111101111111111010111100000100000110001010000111110000000010110100000001111000001111010101011000000000000001000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000001100110111101011010000100001100010010100110000010101011111101101111010110101111010110100000111001100000000111100000001100000000011110000000011011111111100000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000001101011010111101010100000010100010100001010010101010111110111110101101111111111111110111110011000100010000110110000010000000000010010000001110110101011000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000011101011111100110101000100011001001000110100010101010101111101111101110111110101011111100111100110010000001111110000000101111010001000001111011101111101000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000111010101110110101010001000110000100000101000010101010111101111010111010111011111100001111001100010001000000111111000001110000000000000111011101111010110000000000000000000000000000000000000100000000000000000000000000000000000" &
"00000000000000000000000000000000000110101111011011010101000000100010000101010001010010100110111011110101101111111111111110011100111001000100000001111000011000000000000111110110110101111100000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000001110110111101101101010000001101001010010100010101010100111101101011111010111101000011111101111011001100010000111111111110011111111001011011111011110110000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000001110011101011010010100100001010010001101000101001010101010101101101010101010111111100011110011001100010010000011101111100111000000000110110101101101110000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000011010110111101011010010000010100000101010000010101010100101010110101101010011111111111100111001100100010000000000101111111100000000000111111110111011100000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000011101111101010101010010100110000100101000010101010100100101011010101010010111110110111110001100110011001001000000011101101001111110100101010101101111000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000111010101011111010101101000011010010110000010100101001000101010101010101010011111011101111100110011000001000100000000000000111100000000111111110111010000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000110101110110100101000010000100100011001001001010010100010000100000101000000111011010001010110011001001000100000000000001001110000000000010101011101110000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000001110110101110101010011010001101001010100000101001000000000010001000000101001111101011010101011001000100100000010000000000000101111111000111111101011100000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000001101011111101101001010101001010000101000101001000010101000000000001000000011110101101010000101100100110000010000000000000001111110100100010101011110100000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000011110110101010010101101000001001011010000010100010000000001011010000010000011001110110101110010110010010010000000000000010000110000000000011111110111000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000011010111110101000110100100011000010000010101010000001010111111111111101010111101111101100001000110010000000010000010000000110111111101000010101011101000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000011011010101001010101010000010100101100100010001001011111010110111111111101110110101010011010010011001010010000000000000101110111110110100101111010110000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000111101111010100101010101000110001010000010100000101101001010010100101101011110111110110100000011001001000000000010000010110101101000000000011010111100000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000110101101101000101010100001101010100100100000101110010010000000000000010111110110101000101010001101000000000000000011011111110111111110000011011101100000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000001111011101010010010101000011100010100010000011010010010000000101010100001111010001011111010011100100001000001011111101101010111111111111110010110111000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000001110111011000110101000000111101010001000001010101000000000001110110110101110111101101100101000100100100000101100101010111111010110100000000011101101000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000011101010101110110010110000111100010100000101101000100000010100101111001111101101010100011000110110010000010010101011101010101101111011000000010110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000011101111110010110000000011111101000000010110100100001001010100111011011010010110101101101010010010000000001000110010101011110111111110111100101010110000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000111011010101000111000000101111010100000101001000000001010101010111101111101111010101110110010011001001010100100010010101010101101010000000010010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000111011011010100111000000101011000000011011000000100110101011010101001101101010101100111001001001000001111110010001001010101011011111111010000001101100000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000001110111100100101011110000111111100010101100010010001001010101000100111111011111101111100000100101001000010101100100100001000101001111111110000010110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000001111010101010110011101000000101100001010001000000101101101000000001111101011101010000000110110100000000000000001010001010101010101000000001100101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000001101110110101011011110100001110100100100100000100101010010000000111101110110101011011010010010011000000000001111010110000010001011111100000000010011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000011101011001011010101111101001011000010010000010101100000000000011101110011001010101100001001001000000000000100000101111010100101001111111110000011001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000011111101010101111000111110101101100101000010101000000000000001010101011110011011011010101101001000000010110000000000011111000000111010001011001001011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000011010110101111010110011111011110100000001000000000000000000010111101101011010111110100100100100000101101001010100000000101110010011111100000000101001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000001000000000000111110101011010101010001111110101000101000000000000000000001011101010111100111010110010010010000110010110111001010101101001111100011111111110000100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000001000000000000111011010110110110101000001011010100000000000000000000000111111111111110110101011001001010000111010101010001110101001010100001111111000001001000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000001000000000001111110111011011001010000111111001011111111111111110101011100101010010100000010100000101000111010101010101101010100101111010100101111111000000001000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000001100000000000101011011101010100100100111101101010101001010111111010100101010101101011111111011111110111001010101010100101010101010111111010000111111111100000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000001110000000010101010101010101010101010001110101001001101010101111110000000000000010001001001101111011101011010101010101010101010101110101101010110010101011000100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000110000000000010101101101010101001001000011101010010010010100101111111000001010001001010110110101101011001010101010101010101010101101111011100111110000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000111100000000001001010101010110101100000001110100000001010100101011111110100001000100101011011010111011010101010100101001010101001111101110001110111111110000010010000000000000010000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000011110000000000010101010110101101010100000111010101000011010010100111111010000010010010001001101101101001010101010101010101010101011110101101111000100000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000011101010000011000100110101010101010010000011110100101010111100001000111111001000001001101110110010110101010101000101010010101010111011110101111110000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000001111101010100100101010101010100100100100001110010000101010111010010101011110010000010010010011011011000101010110101011010101011101101010011011111111101000001010000100000101000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000111101010111010000100100101010110110000000111101010001010101110100000101111100001000101001100100110011010100010101010010101010111111111011100010101000011000000000001010000101111010000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000011111111010000101010010100110010010010000001110101000101011011011010010111111100010001010010111011001001010101010101001010101101011010011111100000000001110000010000000110010000101010100000000000000000000000000000000000000000000000000000000000000" &
"00000000000000001111111110010100100100100101000100101000001111010010000101011110101000000111100000100101010100101010000101010101010101001001111111101011011111110100000101000000000010001001100010100010101000000000000000000000000000000000000000000000000000000000" &
"00000000000000000001010110100010010010100010100100010101000011101100100010101011110101010101111100000010001010110100110100101010101001010010101010110111100000000000110011101000010100010010010000101111001010010000000000000000000000000000000000000000000000000000" &
"00000000000000000000111100001001001010101000010010001000000001110010010001011101011101000000111110101001010101011000000101001010101010100101111111010111111100000000111000010001000001001000011010000000001100100100000000000000000000000000000000000000000000000000" &
"00000000000000000000000001010100100100101010010001010001000001111101000000100111110111110100010111000000010010100100110010100101010101001010110110100110111111111010110110001000101101000010100110110100100010010000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000010010101010101010100000100100000011111110100010100101111011010001011111010001001010001001000000100101010101001111011011111000101000000111000000010100000011001011001010011011000000010101000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000101001010110101010010000100000011101010000001011011101111111000010111100000100011000010011010101010010010101010110100111110000000001000000000000000100010000001100111001000101001000000100000000000000000000000000000000000000000000" &
"00000000000000000000000000000010000100101001010010101010001000001111011100000100110111011011110000111110000010100000000100010010010010101010111011001101011110101000000000100010001011000101100011000101000000110101010000100000000000000000000000000000000000000000" &
"00000000000000000000000000000000010010101010101011010100100001000111101010000010101010110110111100000111110000010100100010001001101010100101111101011111000101010000000000000001010000101010011000010000101010001000001010000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000100100101001010101101000000000011111010000000010101101101101011010011110000010000001000100101001010101010101101011011110000000000100100000100100100110001000111101011011001100101101000100100000000000000000000000000000000000000" &
"00000000000000000000000000000000010001010100101001010010111010000001110110100001001010110111111111100001011100001000010010001010110101010101111010011101111110101000000000101110000011001100111001100110100110011000000000010000000000000000000000000000000000000000" &
"00000000000000000000000000000001110100001001010110101101010101010000111101010100100101011010101101011100011110000000000000100010010100101011101101011110000101000000000010000000111001001101110010001000111001101110011110100000100000000000000000000000000000000000" &
"00000000000000000000000000000111001110001010100001010110101010101000111111010000010101010101110111110101000111100100001010101001010101010100110100110111100000000001001000101000011000110111001101101010001011100011000000000010010000000000000000000000000000000000" &
"00000000000000000000000000011110101111100001010110101001010100100100001101101000000101010101010101011110100011110000100000010101010101001011101010111011111101010000000010100110100011010100110010010110100100010110001010101000000001000000000000000000000000000000" &
"00000000000000000000000000101011101101000010001001010101010101010101001111010000000100010110101110111011010001111000000001010010101010101010110100111100001011000010101000010001010100101010001010101101111001001000100001010101000000000000000000000000000000000000" &
"00000000000000000000000001111110001100110000100100101010101010101000000111101100000010101010110101101101111010011000001000010100010010010100101010111111000000000000000001010110000111101110101110110011011100101010101101010010101000100000000000000000000000000000" &
"00000000000000000000000110110101100010001000010101010101001010010010100111110010000001010101010110110111101101001010000010001001001000101010110101101011111101010001000000001000111000111011100110011101101110010110010011001001000010001000000000000000000000000000" &
"00000000000000000000001011111010100101010001000010100010101010101010010001101100100010010010011011011101111010100010010000100000101010101001011010111001011110100000011110100111001111011011001001110111010011100011001101100110101010000000000000000000000000000000" &
"00000000000000000000111110100101001000000000001001010101001010010010100011111110001000101001010101101011011111000011000010001010010100010101101001111110000000000101000001111000110110110110010110110101101000011101011100111000000000000000000000000000000000000000" &
"00000000000000000001110111010110010101100010100100100010101010101001000000111010100000000101001010111101101010110000100000100000101010100100110011101111110000000000101010011100101011101101110101001010011111100010100010110001000100101000100000000000000000000000" &
"00000000000000000011010000110101010100010100000001010101010100101010101000111111000000010010101011010110111111011000110000000010010010010011000001110101101111000100000011001010101010111010111111100101101010111100101101000001010001000100000000000000000000000000" &
"00000000000000000111101001011010101010100001000000001001010101010100010000011101010100100100101101011010101011101000010001001001000001011010100011111010000000000010111010110100100101100111010101111011011101101110000000010100001100100000000100000000000000000000" &
"00000000000000001110100101011010000101000100010000101010101010100101100000011110100000000001010010101101110101110110001100000000100100100100000011101111010010000011010101001011111100111011110111011011100110110111101101101011010000010100100000000000000000000000" &
"00000000000000011100110011100100110100000001000000010101010101010101010100001111101001000100101010110110101110110101001000001000010001001010000111110001101000001101010110111110101111001100110110110101011011110111001110010100100101011001000000000000000000000000" &
"00000000000000110111010100011010010000000000000000000101010101001010001000000111010100000010001011010101101111010101000100000010000100010100000110111100000000000010101001010111110011100111101111101010101110101100101001111010111010100000010000000000000000000000" &
"00000000000000111001100111110010000001010101000000000101011010100101010101000111110100000100110010101010111011111011000010000000010010100100000111011111101011001010100101011101111111101111011010001011110101110010101010001011001100001010100100000000000000000000" &
"00000000000010110110100111000100000100100000000000000010101010101010101000000011101001000001001010101101010110101010101001000010000010010000100111100010111000001011111101010110011101011010111100101010011110000000010101110100111101000000100001000000000000000000" &
"00000000000110010011010000001010010010000000000000000001101010101010010101000011111010000010010010100110111011110101010001001000000100001100000111111000000000001110101111101011111111010111101000000100000000001100000010101111000000101010000010000000000000000000" &
"00000000000111011101001010100100010001000100000000100001110101010101101010010001111010000000101010010101011111011010101000100000010001010000001110011111101001011111111011011111011010101101000100110010011001101100110000000000001110101100101000010000000000000000" &
"00000000001111010110101000101010001000000000000000000000011010101010010101000000111010000000000101010101101010110101010100010010000000000100001111100010010000001101101111011110111101010000100110110011001011101101100110011001000010010010010101000010000000000000" &
"00000000011010110100100010101000101001000000001001000000001110110101101010100001111101010001010100101010111011101010111010010000000101010000101011110000000000010111111010110111101000000100101110110011011011101101110110110011000001101010010010000000000000000000" &
"00000000111111011101011010100010000010000000000000000000001111010110101010010000111110100000001001101011010110110010101010001000000000001000001101111111101100011110101111111110110001001101111110111111111111111101110110111011000100010100111001010000000000000000" &
"00000000111100011001000100101000101000000000101000000000000101101010101010100100011101001000010010010101011011011001010101000100000010100000001111001111010000011101111101010101101001101101110111110111011011101111111110111011001000000111000100001100000000000000" &
"00000001101110100011011010010000000010000000000000000000000011111011010101010000011111100010000101001010101101101011011010100100010000000000011111110000000000011011110010101010001101101111111111111011111111111111110111110111011001100000111001010001000000000000" &
"00000001110101010101101001001001001000000100000000000000000001101101011010100000001110110100000010100101010110110101010101000010000101010000001101111101001000000100000100010000000001001000010110111111111011101111101111111110011001000000000000100000010000000000" &
"00000011111101000110010101100000000100000000000000000000000001110101101010010100001111010010001000101001010101101010101010101001000000010000011110010110100000000000000000000000000000000000101111111011011011111011111101110110110011000110000001000000000000000000" &
"00000011011001010011101000000101001000000010000000000000000000111110101010101010000111101010000010010101010101011001010110100001000100000000011111100000000100000000000000000000000000000010110111011111111111101111101111111111111111001100010000011010000100000000" &
"00000101101001101011010101010000000000000000000000000000000000011011101010101001000111111010001001010010101011101010101010101001000000000000011011111110111000000000000000000000000000000101011111111011011011011111011111101101110110011100110001001000100000000000" &
"00001101111011010100100010001010001000010000000000000000000000001110101010100100000111010100000010101001001010101001010101011000100000000000111100111111100000000000000000000000000000010101110111011111111111111111111011011111101110111001100010000100000000000000" &
"00001101110010100111101000010010000000000000000000000000000000001111010101011000100011111011000000000100101010110101001010101010000000000000011111000000000000000000000000000000000001100110110111110111011011010111011111111111101110111001100110000001010000000000" &
"00001001110110110010001011010000001000000000000000000000000000000110110101010010000011101100101010101010010101010010100101101000000000000000010111111010011100000000000000000000000101001010110111011011110111111110111011011011011101110011000100010000000001000000" &
"00011110101011011001001100010101000001000000000000000000000000000111101101001001000001111011000000100100100101101001010101010000000000000000111101111111100000000000000000000000001101001011011111111111011110110110111110111111111111100111011100100001001000000000" &
"00011100100100100100010011001000100000000000000000000000000000000011110101101010010001111101000101010001010110110100101010000000000000000000011101000000000000000000000000000000110100010110110111010110110110111101110111110110111011101110011001100000000000000000" &
"00110110001101110111010100000001000000000000000000000000000000000001111010010100100001110110100000001010001010101001010100000000000000000000111111101000101100000000000000000001011001010101101111110110111110101101101101111111111111011110111001100110000000000000" &
"00111101100111010000001000100110000000000000000000000000000000000001101101101010000001111010100001010001010101010010101000000000000000000000110111111111110000000000000000000110101100010110110110110110101101101111111111111011101110111101110011000100000010000000" &
"00111001010101101101001011010000000000000000000000000000000000000001111010100101010000110110101000001010101010101001000000000000000000000000111100010100000000000000000000001110010000010101011111110111101101011011010111011111111101111011100111001100010000000000" &
"00101110110101100101100110000001000000000000000000000000000000000000111101010010101000111101010001100100010101010100000000000000000000000000011111100001001010000000000000110010101001101110110110110101101011011010110110110111011101110111011110011000100000010000" &
"00111010100111001010010100101000000000000000000000000000000000000000011010101010100000111111001000010010101010110101010101010101010101010100101111111111110000101010101011010100110010101101101110101101011010110110101101110110111011101111011100110001000000000000" &
"01101011110010010101010011000100100100000000000000000000000000000000011111010101001000111010101001001001000101010111111011111111111111101111100001000100101111011010110100001010010010101110110110101101010100101001101111011101110111111101111001110011000010000000" &
"10111010101001001010101001001010000000000000000000000000000000000000011101101010100000011110101000100100101010101010001101010110110101111101110011100000010001010000000000010001001010111011010111101010100101101011011010111011101110111111110111100110000100000000" &
"10111011110101101011010010000000000000000000000000000000000000000000001110111010001000111101010100010010010101010101110110111011011110110110101000110001000101000000100111010101010101101101110101011010101010010110110101110111111101110111101111001100001000000000" &
"01010101110101100101010100010100000000000000000000000000000000000000001110100101010000011110100001010100100101010110101011010101101011011111110100111000010010100001000000000001010101011110011101010010001010101001001011101110111011101110011100111000110000010000" &
"01010110110010110010101010001010100000000000000000000000000000000000000111011010100011111101101001001001010101010101010101011101101110111101011010001100001010100000000000100110000101101011101101000101010101000010010111011011110111111111111101110001100001000000" &
"11010101110101010101100101010000000000000000000000000000000000000000000111101010000101011111010010000100010010101010101010100110110111010111110101001100100001000010001110010101001011011101010010101000000000010101101100110111011111111101110011100011000011000000" &
"01111011010110110000100101001001000000000000000000000000000000000000000011010101000110111010101000100010101000101010101101110101011011111101101110100110001100000000000001000110101011101111011010000000000100100000010011001110111111101111101111001110000100000010" &
"01101010110001101101010100100000000010000000000000000000000000000000000011101010011010101111010000010100010101010100110101011011101101010111111011010011000010001000010010001010001010111010110000100100000000001010001010111011110110111110111100111000011100000100" &
"11111101100110111010010011001000100000000000000000000000000000000000000011110000101101011101001000001001000010000011010101010101111101111010111111101001101001000010000001000100010111010111010010000000000000000000100010101110111101111011110111110001110000010000" &
"01110110110101011001000100110100000000000000000000000000000000000000000011101001111110111110100001000100010101011010010110101110101011011111010101010001000000000010000100010100110110111101100000000000000000000000001100110011110111101111011111000111100001100000" &
"01101101010010110101011001000100010000000000000000000000000000000000000001100111111100111011010100010001001000100101001010110101010110101011111111110100110100000000000000110010101111010110100000000000000000000000000011001111011110111101111100111110000110000000" &
"01110110110101011101001010010001000000000000000000000000000000000000000001101011010110111101000000101000100101010100110101101010101011111110101010101110110000000100011011010000101101101011000000000000000000000000001000111001111011111011110101111000011100000000" &
"10111110110100101010110000001000100010000000000000000000000000000000000001011110111010111101011010000010010010010011010110101010111101001011111111111010001010000000100100010001101101111100000000000000000000000000000010000111010111010111010111100101110000001100" &
"10111010011010011001011110100000010100000000000000000000000000000000000001001011110110111010100000010100100100101010010101010110101011110101001001010101001100000000010111010101011110101010000000000000000000000000000000111010111101111110111110101111100001010000" &
"00111110111111000100101000100100001000000000000000000000000000000000000000110110101101111101010100000010010011010101010101010101111010000000000000000000100100001001001000100001011011011000000000000000000000000000000000000101011111011011110101111100001111010000" &
"00010101000101010010110110100010000000000000000000000000000000000000000011110011111001111010100001010100101000101010101010101111000000000000000000100000000000000001010111010101110101101000000000000000000000000000000000111111101011111110111111100010111000000000" &
"11011100111110101110001010100101010000000000000000000000000000000000000110110101011101110111001000000010001010100101010101110100000000000001000000000010000000010000000110100110111110110010000000000000000000000000000000000000111111010111111100111111110000000110" &
"11011101010111100101010101100100010010100000000000000000000000000000011011010111111011111000100110101000100101010010010110100000000000001000001010100100000000100010111010101011010101010000000000000000000000010000000000001111010101111111100111111110000001011000" &
"10101110101010101001010001100011100100000000000000000000000000000000001111101111110011110111010000000101001000101101101011000010001000010010000000010100010000000000010110100101111110100000000000000000000000000000000000000001011111110100111111101000010111100000" &
"10010101011111101011010100001000000100101010000000000000000000000011101100011010101111101100100001010010010010101010111000000000000000100000000100000000000101010000111111001101110101010000000000000000000000000000000000001010110100101111111010010111111100000000" &
"10111111101101100110011101101000101000100101000000000000000000001011010101101111101111110010000100000001000101010101010000000010000010000000010010101001000000001011010101000111101010100000000000000000000000000000000000000101011111111110101111111101000000000000" &
"01101010110110101011110110010010000010000000010010000000000000001010111111100001001111101101010000010100101011010101000000001000000000100000000010010000001001000101010110001101011110000000000000000000000000000000000000000101101011010111111010010000010001010100" &
"11011111011001100101010101001011010001010000100100101000000111111100101010101110111110110100100010100100101010101110000001000000000010011000101101010000000000100010110110011011101010100000000000000000000010000000000000000010101101101010101111111111111110100000" &
"11100110111010101010110111010100110010100110010011010111111010110111011111101110111111010101001000010010010101010100010000000100010100000111001000100111111110101101011100010101110101000000000000000000000000000000000010000110111111111111111111111111000000000000" &
"11010101111101110101011101010111010010111100101100001010011110111110101010011011111110101001010101001010110101011000000000101000000001111011010110100000000101010010110000011011011010000000000000000000000000000000000000000001010010101010101000000000000000000000" &
"11110111111110011100101011000100101001000011000010011100101010110110010100111011111101100100000010101001010110110000000101000001011111001010101001001111111101010101100100110111011010000000000000000000000000000000000000000111111111111111111111111101110101000000" &
"10110011011010110111010101010010110100001000111010100001001001001010111111001011111010101000101000100101010101000010010000010000100001101110011110100000101011100110000110101101101000000000000000000000000000000000000000000010111110111111111111111111111111111110" &
"01100011111111011101010001011000000101010001001010100101000101101011110111010111110110100101000010010101010110000010000010000001011101010100101010111101011110111000110010111110110100000000000000000000000000000000000000000011101111101010100100100000000000000000" &
"01111100101111000101101100101111010010010100110111010101110010110101111110011111101010010010000101001001011000000000001000101110101011101010110111001001101011000010010110101010101000000000000000000000100000000000000000000110110101111111111111111111010000000000" &
"01101000111011101111101010110010101101101010011000010111010111011011010110111111011010100100010001010101101000010100000010000010101010010011010101111011011010000110011011011110110100000000000000000000000000000000000000000111111111101101001011011111111111000000" &
"01111101001111101010011101011110100100101101000001011001001010101010111101111101101010001001000100101010100001000000101001111010010101101010111110110100101100100011011111011010101000000000000000000000000000000000000000000101010101111111111100000000001010111010" &
"01011111001111100111111010100101110011110101001010100110000101010100010011111101010010100000100101001011000000010100000000001010101010100101000101100011111000110111011110101110100000000000000000000000000000000000000000001111111111010010111111111000000000000000" &
"01011111000011101010111010011111011001011111010101010000111010101011101011101010101001000010001000010101000010100000101110110110101010101001111111011110100100011011111111011010110000000000000000000000000000000000001000000101010111111111100001011111100000000000" &
"00110110011100101011010111010101011000000000110101101011010101011111111010110110100100010000010010101100001000001001010010101101111111111100110101100011010010011011111101011101010000000000000000000000000000000000000000011111111110101010111111000001111100000000" &
"00101110100110101101010101010101111011101100011110110101101011010101011100010101010010001000001010110000100010110100011010111010000001010110101010101110000011011111101110110110100000000000000000000000000000000000000000010111011011111111010101111000000011100000" &
"00101111110101110111101010110100000101110111001011001010011101101011110100000100100001010010101001010001000000011110100000100000011110011000010110110000010011011101111111011010000000000000000000000000000000000000000000011010111111010111111010011111000000001000" &
"00101101110011101101110001011011101010011101100000010101101011001110101000000010001010000010000101100010000101100100001111111111100001101111011000000100010011101111110110111010100000000000000000000000000000000000000000111111110101111100111111000001110000000100" &
"00001111100010111101101110111011010111100110110101101010010100010101110111100000100000101001010101000010000000011101111101101001110101010010110100000010011011101110111111011010000000000000000000000000000000000010000001101011111111011111000111110000011000000000" &
"00001011101101010111111100101110111001011110110110110100101010101010101010111100000001001001001010001000010110110111011111111110010010101011001000010010001001110111111110101101000000000000000000000000000000000000000010111111011111110011111000111100000110000000" &
"00011011101100111101011110110110111001010011101011011011000101111010011011111111000000001010010000001000000110101010110101000111100010001010101010000001001101111110111111110100000000000000000000000000100000000000000011101011110101111101111100001111000011000000" &
"00001011111100001111111011011011110100101100001101010111110111011101011110111011000001010000101000100101001001010101010010110110101011101001001000010001001100110111111010101101000000000000000000000000000000000000001110111110111110010111000111100011100000100000" &
"00000011011100100111101111000110111110101010110101111110101010110111011011011110000000000101000010111011101001111111111101010101010100101010101010001001100110111111111111010100000000100000000000000000000000010000011011111011110101111011100011110000110000010000" &
"00000011111011100001111101010010100010110111010110101011010110101101010111110101010000001000001001001111000111011011101100101101001011101100101000100000100110110111011110110100001000000100000000000000000000000001110111101110011110111100111100111000001000000000" &
"00000010111111100100001111101101010110101110111001011100001011011010111101101101011110000001000011011010010101111110111011011010011100101001101101001000100110111011111110101100000010010000000000001000000000000111011101111011110111011110011100011100001100000000" &
"00000010111011011100010001011111101001101011101101100001100101101101000110110010110111110000011011011100101111010110101010100011100010101101010000000000100110110111111011010000001000000010100100000000000001011101110111011101111011100111100111000110000010000000" &
"00000010111111011100010110110011011110110111011110010111011010110010111001001111101110111101011010110010011101110011111001011100011110101010110010100000110110011111011111101000000001010000101011101001011111110111011111101111011101111011100011000011000010000000" &
"00000010110111111101101011011110111010011100110110101010111101001101101110101010111011111001010101101000101010101011010111010111100101111010100101010000100011011011111110101001001000010010101010101111010101101101111101111011101110011100111001110001100000000000" &
"00000000110110111011100101110111110111001011111110110101101010101111111111001011101101010010101011001011111111111101100001101101101011010001011001000000110110111111111110101000000010010010000101011010111111011111110111011110110111011100111100111000100000000000" &
"00000000101111111111000011011010111101100101010000101111101111101010110101101101101111110100101000101101110101111011011110111011011101101010010011010000100010010111011011010000010000010000110101011011110101111101101101110111111011100111001100011000010000000000" &
"00000000010101111011101001111111101111101010101110010100110111011011011101010101010101001011011111000001011111110110001010111111010111010101110110001000100111011011111110100000000010010010010010101111011111110111111110111111011101110011000110000110010000000000" &
"00000000000101110111011100010101011100101011101011100111011100001101101010010010101101101101110011110111110111011001111101101011110101101001001101100000110010011110111110100000100010010010010010101101101011011111011011011011101110111001110011000110001000000000" &
"00000000001101110111011100000111110111111101011110110001100011110010101101111001010101011110011100110011111101100110000001111110001110001011011001000100000011010111111110100000000000100010110010101101101101111011101111101101110110011101110011100010000000000000" &
"00000000000101110111111001100000111111100111111011011100101110011100110010101111000101100011101101100101011111100001111110110101111001010100110110010000100110110110111101000001000100100110010110110110111101101111111101111110110111001110111001100001000000000000" &
"00000000000101101110111111100100000000011010110111111101010101110111001011011011110110011011011011001111110101101111111101011101010000101011101100100100010110011110111110100100001000100010110010100110110110111101110111110110111011101110011000100001000000000000" &
"00000000000001101111111011101110010001101011101111101110111011011011011101101101011001110110110110010010111110111110101101101010000101001010011001100000000100110111110110000000000001000100100110110110110111110110111110111011011001100110001100010000100000000000" &
"00000000000001001101111111101110011000011111111101011100101101110101100111011011101101011011011001101101101101101011111010111000100100110101110011001000100110101101101110000000010001001100100110010110110110111110110111011111011101110011001100011000000000000000" &
"00000000000000101101110111111100111011000101010111111011110111011111101101010111011010101101110101011011110101111101101011100001010010001001001110010100000100101101111010000000100010001001100110110110110111010110111011011011101100110011000110001000000000000000" &
"00000000000000100101110111011111111011000001011101000100111101110110011011101100110101110011000110101100010110101111111101010110010101001010111001000000100100101011011010000010000010001001100100110110110111011111111111111101101110111001100010001000000000000000" &
"00000000000000001101110111011101110111001100000000101111010111011001101100111011101110101110001111110001111111111010110100100100101000110010100011001010001001101011010100000000000100011001001110100110110111010111011011101101100110011001100011001000000000001000" &
"00000000000000000101100111111101110111011100110000010010101010110010101011001110010011110000001000000011001110110111100001010000010010000101001100110000001001011010110000001000001000010001001100110110110110011011011011101101110110011001110010000000000000000000" &
"00000000000000000100101110011111111111011101110011000101010100000101111101111000101000000011001100011001010111011110010110101101001001001010111010100100000001001110100000000000100000100011001101100110110011011011011011101100110110011100100001000000000000000000" &
"00000000000000000001100110111011101111111101110111100100001000100010001010100010001000110011101110111011111001110101111111111001010010010010100101001000001010010101000000000000000001000110011001101110110110110111011011101110110011001100110001000000000000000000" &
"00000000000000000001000110111011101110111101110111001110011001110010001000100011001101110011101110111101101110101111110110110010101100100101010000100000000010101000000000000010000110000100011001001100110110110111011101101100110110001100110000000000000000000000" &
"00000000000000000000100110111011111110111111111111101110111101110011001100110011001100111011111111011101110111111011011011100100010001001000100111000100000100100000000000001000001000001000110011011101100110110111011001101100110011001100010001000000000000000000" &
"00000000000000000000000100111011011110111011110111101110111001110111011101110111101111111011111111011101110101101101111110101011100010010010101100011000001000000000000000000000010000011001100111011001110110110010011011100110110011001100100000000000000000000000" &
"00000000000000000000000100110011011110111011111111011110111111110111011101111111101110111111101111111111110110110101010101011101110100100101011001100010000001000000000000000000100000100011000110011011101100110111011001101100110110000100000000000000000000000000" &
"00000000000000000000000100110011011101111111101111111111111011110111011101110111111111111011111111011111110011111011101011101111100011001000010011000100000010000000000000000000000011000010001100110011001101110110011011101100110010001000100000000000000000000000" &
"00000000000000000000000010010011011101110111111111011110111111111111011110111111101110111111111111111110111101010110101101101101001000010010100100011000000000000000000000000000000100001100011000110011001100100100110011001100110010001000000000000000000000000000" &
"00000000000000000000000000110011001101110111011111011111111011110111111111111011111111111111111111011111111110111101111101111010100101100101001001100010000000000000000000000000000000010000110001100111011001100110110011001000110010001000000000000000000000000000" &
"00000000000000000000000000010010011101110111101111111101111111111111011101111111101111111111101111111110110110010111110100001010100100010010010010001000000000000000000000000000000001000001100011001110011001101100110010001100100010000000000000000000000000000000" &
"00000000000000000000000000000010011001110111011110111111111011110111111111111011111110111011111111011110111111101110101111111111111110100100100101110001000000000000000000000000000000000110000110011100110011001000100011001000100010000000000000000000000000000000" &
"00000000000000000000000000000010001101100111011110111101111111111111011111111111101111111111110111111110111011101011110101010101010110001000001000100010000000000000000000000000000000001000000100011000100011001001100110011001000000000000000000000000000000000000" &
"00000000000000000000000000000001001000100111001110111101111011101111111110111011111111111011101111011110111111100111001010110110111100110011001011001100000000000000000000000000000000000000011000110001000110010001000100000001000000000000000000000000000000000000" &
"00000000000000000000000000000000001001100111011100111011111011111111011111111111101110111101111111101110110111101101111101011111111010000100010010010001000000000000000000000000000000000000100001100011001100010010000100010000000000000000000000000000000000000000" &
"00000000000000000000000000000000001000110110011100111001110111101111011101111011111111111111110111011110111111101010101101101010101011011000100100100110000000000000000000000000000000000000000010000100001000100010001000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000001100011001100111011110111101110111111111111101110111011101111011101110111001110111010101010010101111001001001001001010000000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000010011100111001110111101111111101110111101110111011101111011101110111011110101101101101110110111010010010010110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000100010011000110011110111001110111111110111011110111011101111011101110111011100001011010111010011100000100100101100101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000010001000110011100111011110111101110111011110111001101110011101100111001101110110111101110101010011001000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000010011000110011100111001100111001100111001100111011100110111001100110011101110011010110100100000100010010100110110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000110011000110011101111011100111011101110011001110011001101110011001100001111011011011111111000100010001001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000001000100011000110011100111011101110011100110011101100111001100100110001100110001101011101101100001001001010110100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000100010001100011001110011001110011001110011001100110011001100110011001000000111101101110101111000010100101101001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000010000100011001110011001100011000100110001100110011001000100110000000000001111011011000011100100001010011010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000001000110001100010001100110001100110011001100110001001000000000000000000010111100101101001010010011101110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000001000100011000110001000110011000100010001000100010001000000000000000000001100010111010010000100101011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000100010000100011000100001001100110001000100000000000000000000000000000001101101010100101001010110011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000001000010001000010001000000010000000001010000000000000000000000000010101011111010010111011100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000010000010000100000000000000000000000000000000011101011100101000100100000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111011001000001000000000000000000000000000000000111111010010110111010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111101100010100000000000000000000000000000000000101011001100001000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000010000000000000000000000000000000000000000001110100001000000000000000000000000000000000000000011110010011010011110001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000001111110000000000000000000000000000010000000011110100000000000000000000000000000000000000000000001000100000101101000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000011011110000000000000011110000000000111100000011011010100100000000000000000000000000000000000000001011011010010010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000111001011000000000000111011100000001111110000111010010000000000010111000000000000000001000000000001110111000101011000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000111010110000000000001110001010000001101010000111100100010100000010111000000000000000011111000000001011101100001010110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000110000001100000000000101001111000011010001001111010001000000000101011100000000000000111011110000001101010110101111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000101000010010000000001101100000000011100011011010100100001000001101110110000000000001111101010000001011111110010000100000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000111001100100000000001010100101000111100001001101100000100000011100110001000000000001111001111000001100010000001110000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000110100110100000000000000011000100111011100011110001000000000011001011001000000000001111000001000001111000011101001000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000011000110010000000000100000101000111010110111101000010100000111000110001000000000001111000000000001110110000011100000011110111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000010100011000000111111111100000100100010101101010100001000000111100101001000101100001111011010110001110100101000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000011010010000001111101111110000100110001001110100010100000000110110001101011111100001110111110000011011010010110000000101111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000011100011000111111011010111100000000000111110101000000000000111110001010111000100011110001011010011010101000000000000111101111001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000001010001000111101101101111111110100001101011000000010000000111010001101001010010000100001011000011100100011000000000101101110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000010000010100001001110000100010100011010111011101110100001000000000101101001011011101000000110001010100111010011000000000001111001000111000000100000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000001011101101001110001001101000001010001001110111111010011001000001101000110110000101011110001000010000101010011111000010100001001011010001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000101010001000000000000101000000100001011111101110110100101000010001011000101001001011001010010100101000001000111010001000100000011110010010111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000001011110101010001010010010101000001110111010101101001001100100000000010000101100000100001110001110001100010101011010100101111000010100110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000011111111101000000001111101111011111101110111001000000011110001000011000100100101000100010110000100010010000010101110000000101000101110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000011111111100001000111111101110111010101100000100101000101000010000001100000000000000000000001001011000100000101110000101000011000011000100011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000001111111110100001111110111001101011000010101000000011110101000010010111100000000000011000000000101000010000011101010000010010100101101101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000111111011010011110010101101110000101000000001000111101000100001000100111110111011111100100000011000001000001101000010011001110010011000011000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000011010001010111001000010100001010000000100000011100100010000000000100010111011110111111111100001000010000011011010000010001010010010001010001011111111000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000010100000111000000010010100000001000000000111110101000000000100001011001101011010110111111000000000000110101000000101000101001010000001111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000010100001100001010010000000010000010010001010100000000000000000000000010101010111011111111001000000100111010100000100011000000100000110101011111111100000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000001000100111001001000000000001010100111101010010000000000000001001001000101001010001111100100000001111000001001000111111000100010111010111111010100000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000001100000100000001000000001000001011010100000001011000100000000010001010010100000001110100000001110110000000101111011100000101100100010100001000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000011110000000000000001000000100000001011000000011101000010001100100010111000000000000000001010000001110000001001011010000001001111000110000010001001101001111000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000111111100000000010111111110000000000000100001111010101000001010001010111110000000001001000000111110010100100011101100100001001111110001100000100110110001010000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000111110101000101000010111011000011010000001110110100100000000100111110011111101000000000001000100010010000010011101010000000100111111111101000010011011010110000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000111111000011111111001001101111111111110011111001010000000001000110111001011101101010000000001001101010100100111100000001010001111011111011100001010110011100000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000101110010111111111100100010000000000000111101001000010001000000111101000100100110111010000001100111010010000111111010100010000111101011101110001011110010100000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000101010000011111111101101101011010000100101110100001000011110001111111010100001100010001000111100011000010001011010100000001001111000101011110001101000101000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000001010010100111111111010010010100101110000111010000100000111111000111110101111000111001001011111110101100010001101101001000000000111001011101111000100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000001100001100001111111000000100001010010011111010110000001001010101111011101010100011000001100111110010110010001110010100000100100111100010101111001000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000110101010100001000000000000100000000011110000000000000010101101111111010101100101100010101111100001011000011111000000000010101110100001001111000010100010000000000000100000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000101000100001001010111010000110000000111100000000000011001000100101111101010010010100001001111111000100001001101110000100110100001110001011011100010000000000000000010000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000010100111000101010000100001111010100111000001000001101100010110010001000001000000110001011111001100100000001110101010000110000000011000001111100100000000000010000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000011000010100000101010000011101100000111000100100010101010101010011110101000000000001000111110010110010010011011010000000101000110011100010010110000000000001100000000001010101000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000001100001100100000000010011110011100111000000000101101000111110101011000000011111100000101010010010000000011101101000001010100001000100000111110000010000111111000101010010101100000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000110001010000100000000111101000100110000000000110101010001010000100110001111111111000011011001010010001011110010100000100000001100110000010110001000001101111000000101010101110000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000010100110010001000000111111110000110011010011010101001111001000101000011111111111001000101010010010000110111000000001101000010100001100101011000100011110111100001001010111111100000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000010100011000100000001111001110110110001011010101010000010010000010000111101111110111100000000000000001101011010000000110100000111000111001101000000111101111110001011011000111110000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000001000010100000100001111101011001011010000000010100101101011000000001110010000101111110101000000010111110101000000000110110000010100111000101101010111101101110010101000000001111100000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000001101001000100000011110011101101011000101101000100000100011000100001000000000011101011101010010101101010111010000010010011000101010011000101100001111101011111000000000000100111110000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000100000110001010001010100110100100101110111010000010010101010000011010100000110101010010111111111100101001100000010110000001001000101100101010011111000110111000001100010011000010000000100000000000000000000000000000000000000000000" &
"00000000000000000000000000000000010000100000000001100010010110100001111011111110000100011000101001010001010001000011111110111011010101110000100001000100000000110001100001010101110011001111100000000001101001000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000111110000000010000010001011010101010100011110101011111100000110000100001010110000000111111011101101001010001101000000010101110000000000000110000010001010001111010000000000001010001010100000000000000000000000000000000000000000000000000" &
"00000000000000000000000011111111110000001000000101110001001011010011111010110101110000110000000100000000101011110110010100110010100011010000000000011011110100000000000000000001010010111101100010101001110101100000000000000000000000000000000000000000000000000000" &
"00000000000000000000000111111110011111000000000000101000101010010111111101010110100001100000000000011111111111001101010100001000000110101001000001001001111111110111100000000000100001011100000001010110000110000000000000000000000000000000000000000000000000000000" &
"00000000000000000000001111111110001011111010001000111100100101010001111100101011111001001010010000111110110101100100010001000000001110010000000000000010100111111111111111111000000010101010110100101001101000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000001111111101000000011110100000110100000010010001111100010100010100100100001110110101110100010010000000000000111011000100000000000100101010011101111111111110000101111001000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000011101011010100000101110100111101000100010001111111000001011010000001011111111001010101000000000000000001110101000000000000000000000110101100111011111111000000010101100000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000100100011101001000000011010101010001110011001111011100000101010000000111110101101001000000000000000100011101000000000000000000000100001001101101111110111100001010010110000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000001010011011010101000000010111110000110001000111101111000001001000001111101110101010001000000010010001111010101000001011010010000001000010010101000000001110000100010010000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000100101001110110100010000000010101010010010100110010011011000100001011110000001000000000000001100000111100101000000011100010000000000001000001010100000000000000000101100000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000010010000011111010101000000011010001011001010101001001000110010100011100000000000000000001110010001111110010000000011000010011010000000001000010001111111110100000010110000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000010110000010111010010000011101000101000000010000100100101001010011000101001000000000010001000111001001000000010010110010000000101000000010100010101111111111000010010000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000001011101000001010101000001011000011001100011110001000100010100011001110100000000100000100001110100100000001010010011100000100001010000000000010101111111111110101100000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000010101001000001010010011101001011000000001101100010010000010011001111000000000110000000110111110101000011010010010010000000101011100000000010011111111111110010100000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000010110010000001000001111000101001101010111010001001001010100011110100000010001000011111010100000001000010010010101010010111010111001011000011111111001100010000000000000000000000000000000100000000000000000000000000000000000000000" &
"00000000000000000000000000000000000001010010000001010101100010100100010110101000110000001000011101011101100010100111110101010100010001101010010011000101111011011000010101111111101010100101000000000100000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000001100100010001111000101000001100010100100101000100000111101010010110100000011011100010000010101101011010010001001111101101010101011011111010101001010000001011111000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000001001110001010100000100011000010101000010100000100011100101010010001011110110010100000001000100010010011010011111100010100010101011100110110000110001011111111000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000011000101101100010100110100001100000001010000000111001001010100100111111010100000001000010010101001010000010111110101000100101001011011010010100010111110000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000110000010110100000011101000000110101001101000000111000100000001001111000001000100010001000110010010010011010111100001000001000011010101100001010001101001101100000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000001100010101011010000111010101000100100000010000100101000001001010001110100001000000000001000001011010011001001001101010100000010101101101000101000101111010011000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000111000101010101000001111101010010011001000011010000111100000101000011100000000001001010101100010010000101010110110001000000000000101010111000010000011000011010000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000001010001010100110100001111010000010000000000001000000101010010110100111100000100100001000000100001010010010001010101001100110010111011101100001001000100000100010000000000000000100000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000001100010101000000000001111001101010010110100001010000101111000010100111000000000000110110001011000010110011010101010010101000000011110110100100010000010100101100000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000001110101110000100101001110010101000100000000000100100110010101011100111000010000000110010100100100001000001001010110001010100011000101000000000100101000000010000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000010010111101111001000011100101000111110010000010100000010000010101000001000110000000000001110000000010010010010010001100100100101100100010000010001000100000000101100000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000011011101001110010100010111111000010001000100000000000000001000010101000101100110001000101011101000000010101000000011000100110001010100001000000100010000000001011010000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000001101000100111010101001001111111000001000010001001000010000000001100100100010010011000000111111100010100000100100010001001010000010101000010101010000000001001010100000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000110001010101010101101001001111110000100000000100000001000000000111100010000000000011001100001111010101001000010010010010000101010010100100000010101000000000001000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000100101010010001101110100011111101010000101000000000000000100001111100000000010101001001010000011101000100000010100000001000101000001000100101000001011100010010000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000001111010101000110101000011111101010110100101001010000001000111111000000010000110100100000000100110111001000000010000001000101000100011000010101000010110000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000001111101100000000000000001010100011011011010100100100100000001111100101110000000110010000101000010010100110100000100100000000010100000010100000101010100010100000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000011101111000010100001001000010100011111101101010101001000000011111010111111100001110100000000000000001110100100100001000010000010101010010110010001011111110010000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000001110101101101010100010100001101010101011111111010100010011111100001111100010101100000010010010001000110101001000000001000000010100101001010000000111111110011000000000000000000000000000000010000000000000000000000000000000000000000000000" &
"00000000000000000000000000101110110010000001000100010100000000000000000101011000111111000001000011101001100000111101101010110011010100010010000000000001011101000010000001011111111001100000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000011001000010000100010101001110010100010000100000000011111100000010010100101010101000101010000000001001101010011111111101001001011111000100001001111111111100100000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000100101000100001000000000011010101000100000000000111111000000001000010010101010100100101000000000100110101001011111111110000111111101010000100111111111100100000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000010101001000000000100000000010101011001000100001111100000000100101000000001010100001000000000000000111010100101101101000000111111100100000010001111111101010000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000100100010100000000000000001001000100100001011110000000010001010000000001111010000000010100000010001100010010111000000000111111100100001000000111110101100000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000010010000000000000000000000000000000000100011100000001000100101110100001101101110111010010000000001000100010010000010100111111100100000101000010000110000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000011011101000000110000000100101000110010010000101101001000100100100010100000010011011010101010000000000100000100101000100101000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000010010001000001100001010010100000011001010000100010110110101000000010010000000000101001010110011000000100000000010111101100000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000111101010000000000010001010000000001101001010011011010101000100000011010100000010000110111100001111110000000000000010101000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000111101010000010001001010100010000000010100000011110101001010101010000101010101000100001101000000000101100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000111011100000011101010110101010101000000011010000001010100100000000000000100000001101000110010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000011101100000010011011100100100100010001000010000000000000000001010100000001010001110110000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000001110000000010001101010101010010101010000000100000000100010000110010001000000101110000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000001000000000001000001011010101001101001110000001000000010100010100100000100000000001000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000101010000101011000000111100000110000000001010100011001010000111000000000000000100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000010101010011100000010010110000000000000010101000011001010010001000000001010001010000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000011101000000100000001101001000000000000010101001010000100010001000000000001000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000011110111000000000001010001011101000000101010001110000110110100000000000010000001111010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000001010000000000000000100100110101000001110100000100000010010100000000000000110001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000111010100001111010000000000110011010000000000000001011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100011111100000111010101000000011001100000000000000010100011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101101100000110101000000000001001010000000000000000010101100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000111000000011110100000000001001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000010110000000000001100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011010000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" &
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

  SIGNAL dmem : std_logic;
  
BEGIN


  ----------------------------------------------------------------
  hps : hps_io
    GENERIC MAP (
      STRLEN => CONF_STR'length)
    PORT MAP (
      clk_sys            => clksys,
      hps_bus            => hps_bus,
      conf_str           => to_slv(CONF_STR),
      buttons            => OPEN,
      forced_scandoubler => OPEN,
      joystick_0         => OPEN,
      joystick_1         => OPEN,
      joystick_2         => OPEN,
      joystick_3         => OPEN,
      joystick_4         => OPEN,
      joystick_5         => OPEN,
      joystick_analog_0  => OPEN,
      joystick_analog_1  => OPEN,
      joystick_analog_2  => OPEN,
      joystick_analog_3  => OPEN,
      joystick_analog_4  => OPEN,
      joystick_analog_5  => OPEN,
      buttons            => OPEN,
      forced_scandoubler => OPEN,
      status             => status,
      status_in          => status_in,
      status_set         => status_set,
      status_menumask    => status_menumask,
      new_vmode          => new_vmode,
      img_mounted        => OPEN,
      img_readonly       => OPEN,
      img_size           => OPEN,
      sd_lba             => std_logic_vector'(x"0000_0000"),
      sd_rd              => '0',
      sd_wr              => '0',
      sd_ack             => OPEN,
      sd_conf            => '0',
      sd_ack_conf        => OPEN,
      sd_buff_addr       => OPEN,
      sd_buff_dout       => OPEN,
      sd_buff_din        => std_logic_vector'(x"00"),
      sd_buff_wr         => OPEN,
      ioctl_download     => OPEN,
      ioctl_index        => OPEN,
      ioctl_wr           => OPEN,
      ioctl_addr         => OPEN,
      ioctl_dout         => OPEN,
      ioctl_wait         => ioctl_wait,
      rtc                => OPEN,
      timestamp          => OPEN,
      uart_mode          => std_logic_vector'(x"0000"),
      ps2_kbd_clk_out    => OPEN,
      ps2_kbd_data_out   => OPEN,
      ps2_kbd_clk_in     => '1',
      ps2_kbd_data_in    => '1',
      ps2_kbd_led_use    => std_logic_vector'("000"),
      ps2_kbd_led_status => std_logic_vector'("000"),
      ps2_mouse_clk_out  => OPEN,
      ps2_mouse_data_out => OPEN,
      ps2_mouse_clk_in   => '1',
      ps2_mouse_data_in  => '1',
      ps2_key            => ps2_key,
      ps2_mouse          => OPEN,
      ps2_mouse_ext      => OPEN);
  
  sconf<=status(8 DOWNTO 4);
  vga_sl<="00";
  
  ----------------------------------------------------------
  --ipll : pll
  --  PORT MAP (
  --    refclk   => clk_50m,
  --    rst      => '0',
  --    outclk_0 => clksys,
  --    outclk_1 => clksys2,
  --    locked   => pll_locked
  --    );
  clksys<=clk_50m;
  ----------------------------------------------------------
  VideoGen:PROCESS (clksys) IS
  BEGIN
    IF rising_edge(clksys) THEN
      calt<=calt+1;
      IF calt=7 THEN calt<=0; END IF;
      
      IF calt=0 THEN
        gce<='1';
      ELSE
        gce<='0';
      END IF;
      
      IF gce='1' THEN
        IF ghcpt<ghtotal-1 THEN
          ghcpt<=ghcpt+1;
        ELSE
          ghcpt<=0;
          IF gvcpt<gvtotal-1 THEN
            gvcpt<=gvcpt+1;
          ELSE
            gvcpt<=0;
            gfl<=gfl XOR inter;
          END IF;
        END IF;
        
        gde<=to_std_logic(ghcpt<ghdisp AND gvcpt<gvdisp);
        ghs<=to_std_logic(ghcpt>=ghsyncstart AND ghcpt<ghsyncend);
        gvs<=to_std_logic(gvcpt>=gvsyncstart AND gvcpt<gvsyncend);
      END IF;
    END IF;
  END PROCESS;
  
  ----------------------------------------------------------
  -- MIRE
  MireZ:PROCESS (clksys) IS
    VARIABLE t : std_logic;
    VARIABLE d : unsigned(8 DOWNTO 0); -- RRRGGGBBB
    VARIABLE ghcpt_v,gvcpt_v : natural RANGE 0 TO 4095;
    VARIABLE ghdisp_v,gvdisp_v : natural RANGE 0 TO 4095;
    
  BEGIN
    IF rising_edge(clksys) THEN
      IF gce='1' THEN
        IF double='1' THEN
          ghcpt_v:=ghcpt / 2;
          gvcpt_v:=gvcpt / 2;
          ghdisp_v:=ghdisp / 2;
          gvdisp_v:=gvdisp / 2;
        ELSE
          ghcpt_v:=ghcpt;
          gvcpt_v:=gvcpt;
          ghdisp_v:=ghdisp;
          gvdisp_v:=gvdisp;
        END IF;

        --dmem<=dragon(ghcpt + gvcpt * 260);
        
        CASE mire IS
          WHEN 0 =>
            t:=test(
              (ghcpt_v + gvcpt_v * 320)
--pragma synthesis_off
              MOD (320*128)
--pragma synthesis_on
              );
          WHEN 1 => -- Cadres
            t:=to_std_logic((ghcpt_v=0 OR ghcpt_v=ghdisp_v-1 OR
                             gvcpt_v=0 OR gvcpt_v=gvdisp_v-1) AND
                            ghcpt_v<ghdisp_v AND gvcpt_v<gvdisp_v);
            t:=t OR to_std_logic((ghcpt_v=32 OR ghcpt_v=ghdisp_v-33 OR
                                  gvcpt_v=32 OR gvcpt_v=gvdisp_v-33) AND
                                 ghcpt_v<ghdisp_v AND gvcpt_v<gvdisp_v);
            t:=t OR to_std_logic((ghcpt_v=64 OR ghcpt_v=ghdisp_v-65 OR
                                  gvcpt_v=64 OR gvcpt_v=gvdisp_v-65) AND
                                 ghcpt_v<ghdisp_v AND gvcpt_v<gvdisp_v);
            t:=t OR to_std_logic((ghcpt_v=96 OR ghcpt_v=ghdisp_v-97 OR
                                  gvcpt_v=96 OR gvcpt_v=gvdisp_v-97) AND
                                 ghcpt_v<ghdisp_v AND gvcpt_v<gvdisp_v);
          WHEN 2 => -- Cadrillage
            t:=to_std_logic((ghcpt_v MOD 16)=0 AND (gvcpt_v MOD 16)=0);
            
          WHEN 3 => -- Lignes diagonales
            t:=to_std_logic((ghcpt_v+gvcpt_v) MOD 16 = 0);
            
          WHEN 4 => -- Bandes diagonales
            t:=to_std_logic(((ghcpt_v+gvcpt_v)/16) MOD 2 = 0);
            
          WHEN 5 => -- Damier
            t:=to_std_logic((ghcpt_v/16) MOD 2 = (gvcpt_v/16) MOD 2);
            
          WHEN 6 => -- Cadrillage fin
            t:=to_std_logic((ghcpt_v MOD 4)=0 AND (gvcpt_v MOD 4)=0);
            
          WHEN 7 =>  -- Lignes Horizontales fines 
            t:=to_std_logic(ghcpt_v MOD 2=0);
            
          WHEN 8 => -- Lignes verticales fines
            t:=to_std_logic(gvcpt_v MOD 2=0);

          WHEN 9 => -- Cadrillage diagonal
            t:=to_std_logic((ghcpt_v+gvcpt_v) MOD 16 = 0) OR
                to_std_logic((ghcpt_v-gvcpt_v) MOD 16 = 0);
            
          WHEN 10=> -- Damier diagonal
            t:=to_std_logic(((ghcpt_v+gvcpt_v)/16) MOD 2 = 0) XOR
                to_std_logic(((ghcpt_v-gvcpt_v)/16) MOD 2 = 0);
            
          WHEN 11 =>
            t:=to_std_logic(((ghcpt_v+gvcpt_v)/8) MOD 2 = 0) XOR
                to_std_logic(((ghcpt_v-gvcpt_v)/8) MOD 2 = 0);
            
          WHEN 12 =>
            t:=to_std_logic(((ghcpt_v+gvcpt_v)/128) MOD 2 = 0) XOR
                to_std_logic(((ghcpt_v-gvcpt_v)/128) MOD 2 = 0);
            
          WHEN 13=> -- 
            t:=to_std_logic((ghcpt_v MOD 32)=0 AND (gvcpt_v MOD 32)=0);
            
          WHEN 14 =>
            t:=dragon((ghcpt_v + gvcpt_v * 260)
--pragma synthesis_off
                      MOD (260*400)
--pragma synthesis_on
                      );
            
          WHEN 15 =>
            t:=NOT dragon((ghcpt_v + gvcpt_v * 260)
--pragma synthesis_off
                          MOD (260*400)
--pragma synthesis_on
                          );
        END CASE;
        t:=t OR to_std_logic((ghcpt_v=0 OR ghcpt_v=ghdisp_v-1 OR
                              gvcpt_v=0 OR gvcpt_v=gvdisp_v-1) AND
                             ghcpt_v<ghdisp_v AND gvcpt_v<gvdisp_v);
        
        ----------------------------------
        gr<=(OTHERS =>t);
        gg<=(OTHERS =>t);
        gb<=(OTHERS =>t);
      END IF;
    END IF;
  END PROCESS;
  
  ----------------------------------------------------------
  KeyCodes:PROCESS (clksys,reset_na) IS
  BEGIN
    IF reset_na='0' THEN
      NULL;
    ELSIF rising_edge(clksys) THEN
      key_0<='0';      key_1<='0';
      key_2<='0';      key_3<='0';
      key_4<='0';      key_5<='0';
      key_6<='0';      key_7<='0';
      key_8<='0';      key_9<='0';
      key_q<='0';      key_w<='0';
      key_e<='0';      key_r<='0';
      key_t<='0';      key_y<='0';
      key_u<='0';      key_i<='0';
      key_o<='0';      key_p<='0';
      key_a<='0';      key_s<='0';
      key_d<='0';      key_f<='0';
      key_g<='0';      key_h<='0';
      key_j<='0';      key_k<='0';
      key_l<='0';      key_z<='0';
      key_x<='0';      key_c<='0';
      key_v<='0';      key_b<='0';
      key_n<='0';      key_m<='0';
      key_space<='0'; 
      key_return<='0';
      
      --------------------------
      ps2_key_delay<=ps2_key;
      IF ps2_key_delay(10)/=ps2_key(10) THEN
        CASE ps2_key(7 DOWNTO 0) IS
          WHEN x"45" => key_0<=ps2_key(9);
          WHEN x"16" => key_1<=ps2_key(9);
          WHEN x"1E" => key_2<=ps2_key(9);
          WHEN x"26" => key_3<=ps2_key(9);
          WHEN x"25" => key_4<=ps2_key(9);
          WHEN x"2E" => key_5<=ps2_key(9);
          WHEN x"36" => key_6<=ps2_key(9);
          WHEN x"3D" => key_7<=ps2_key(9);
          WHEN x"3E" => key_8<=ps2_key(9);
          WHEN x"46" => key_9<=ps2_key(9);

          WHEN x"15" => key_q<=ps2_key(9);
          WHEN x"1D" => key_w<=ps2_key(9);
          WHEN x"24" => key_e<=ps2_key(9);
          WHEN x"2D" => key_r<=ps2_key(9);
          WHEN x"2C" => key_t<=ps2_key(9);
          WHEN x"35" => key_y<=ps2_key(9);
          WHEN x"3C" => key_u<=ps2_key(9);
          WHEN x"43" => key_i<=ps2_key(9);
          WHEN x"44" => key_o<=ps2_key(9);
          WHEN x"4D" => key_p<=ps2_key(9);

          WHEN x"1C" => key_a<=ps2_key(9);
          WHEN x"1B" => key_s<=ps2_key(9);
          WHEN x"23" => key_d<=ps2_key(9);
          WHEN x"2B" => key_f<=ps2_key(9);
          WHEN x"34" => key_g<=ps2_key(9);
          WHEN x"33" => key_h<=ps2_key(9);
          WHEN x"3B" => key_j<=ps2_key(9);
          WHEN x"42" => key_k<=ps2_key(9);
          WHEN x"4B" => key_l<=ps2_key(9);
                        
          WHEN x"1A" => key_z<=ps2_key(9);
          WHEN x"22" => key_x<=ps2_key(9);
          WHEN x"21" => key_c<=ps2_key(9);
          WHEN x"2A" => key_v<=ps2_key(9);
          WHEN x"32" => key_b<=ps2_key(9);
          WHEN x"31" => key_n<=ps2_key(9);
          WHEN x"3A" => key_m<=ps2_key(9);
                        
          WHEN x"29" => key_space<=ps2_key(9); -- SPACE
          WHEN x"5A" => key_return<=ps2_key(9); -- RETURN
          WHEN OTHERS => NULL;
        END CASE;
      END IF;
    END IF;
  END PROCESS KeyCodes;

  ----------------------------------------------------------
  Keys:PROCESS(clksys) IS
  BEGIN
    IF rising_edge(clksys) THEN
      IF clkdiv < 10_000_000 THEN
        clkdiv<=clkdiv+1;
      ELSE
        clkdiv<=0;
      END IF;
      
      IF key_a='1' THEN iauto_n_i <=NOT iauto_n_i; END IF;
      IF key_b='1' THEN sel<=0; END IF;
      IF key_c='1' THEN sel<=1; END IF;
      IF key_d='1' THEN sel<=2; END IF;
      IF key_e='1' THEN sel<=3; END IF;
      IF key_f='1' THEN oauto_n_i <=NOT oauto_n_i; END IF;
      IF key_g='1' THEN sel<=4; END IF;
      IF key_h='1' THEN sel<=5; END IF;
      IF key_i='1' THEN sel<=6; END IF;
      IF key_j='1' THEN sel<=7; END IF;
      IF key_k='1' THEN mire<=(mire +1) MOD 16; END IF;
      IF key_l='1' THEN
        iauto_n_i<='0';
        oauto_n_i<='0';
        himin_i<=0;
        himax_i<=ghdisp-1;
        vimax_i<=0;
        vimax_i<=gvdisp-1;
        move<='0';
      END IF;

      IF key_m='1' THEN double<=NOT double; END IF;
      IF key_n='1' THEN inter<=NOT inter; END IF;

      inc<='0';
      dec<='0';
      
      IF key_o='1' THEN
        inc<='1';
        delta<=1;
      END IF;
      IF key_p='1' THEN
        dec<='1';
        delta<=1;
      END IF;
      IF key_9='1' THEN
        inc<='1';
        delta<=10;
      END IF;
      IF key_0='1' THEN
        dec<='1';
        delta<=10;
      END IF;

      IF key_1='1' THEN
        move<=NOT move;
        dir<='0';
      END IF;
      IF key_2='1' THEN
        move<=NOT move;
        dir<='1';
      END IF;

      IF move='1' AND dir='1' AND clkdiv=0 THEN
        dec<='1';
      ELSIF move='1' AND dir='0' AND clkdiv=0 THEN
        inc<='1';
      END IF;
      
      
      CASE sel IS
        WHEN 0 => IF inc='1' THEN himin_i<=himin_i+delta; ELSIF dec='1' AND himin_i>=delta THEN himin_i<=himin_i-delta;  END IF;
        WHEN 1 => IF inc='1' THEN himax_i<=himax_i+delta; ELSIF dec='1' AND himax_i>=delta THEN himax_i<=himax_i-delta;  END IF;
        WHEN 2 => IF inc='1' THEN vimin_i<=vimin_i+delta; ELSIF dec='1' AND vimin_i>=delta THEN vimin_i<=vimin_i-delta;  END IF;
        WHEN 3 => IF inc='1' THEN vimax_i<=vimax_i+delta; ELSIF dec='1' AND vimax_i>=delta THEN vimax_i<=vimax_i-delta;  END IF;
        WHEN 4 => IF inc='1' THEN hmin_i <=hmin_i+delta;  ELSIF dec='1' AND hmin_i>=delta THEN hmin_i <=hmin_i-delta;  END IF;
        WHEN 5 => IF inc='1' THEN hmax_i <=hmax_i+delta;  ELSIF dec='1' AND hmax_i>=delta THEN hmax_i <=hmax_i-delta;  END IF;
        WHEN 6 => IF inc='1' THEN vmin_i <=vmin_i+delta;  ELSIF dec='1' AND vmin_i>=delta THEN vmin_i <=vmin_i-delta;  END IF;
        WHEN 7 => IF inc='1' THEN vmax_i <=vmax_i+delta;  ELSIF dec='1' AND vmax_i>=delta THEN vmax_i <=vmax_i-delta;  END IF;
        WHEN OTHERS => NULL;
      END CASE;

      IF oauto_n_i='0' THEN
        hmin_i<=0;
        hmax_i<=hdisp-1;
        vmin_i<=0;
        vmax_i<=vdisp-1;
      END IF;
    END IF;
  END PROCESS Keys;

  himin<=himin_i;
  himax<=himax_i;
  vimin<=vimin_i;
  vimax<=vimax_i;
  hmin<=hmin_i;
  hmax<=hmax_i;
  vmin<=vmin_i;
  vmax<=vmax_i;
  iauto<=NOT iauto_n_i;
  
  ----------------------------------------------------------
  i_ovo: ENTITY work.ovo
    PORT MAP (
      i_r     => gr,
      i_g     => gg,
      i_b     => gb,
      i_hs    => ghs,
      i_vs    => gvs,
      i_de    => gde,
      i_en    => gce,
      i_clk   => clksys,
      o_r     => vga_r_u,
      o_g     => vga_g_u,
      o_b     => vga_b_u,
      o_hs    => vga_hs,
      o_vs    => vga_vs,
      o_de    => vga_de,
      ena     => ovo_ena,
      in0     => ovo_in0,
      in1     => ovo_in1);

  vga_r<=std_logic_vector(vga_r_u);
  vga_g<=std_logic_vector(vga_g_u);
  vga_b<=std_logic_vector(vga_b_u);

  vga_f1<=gfl;

  ce_pixel<=gce;
  
  clk_video<=clksys;
  
  audio_l<=x"0000";
  audio_r<=x"0000";
  audio_s<='1';
  audio_mix<="11";
  
  ovo_in0<=
    CC(' ') & -- 1
    CN(to_unsigned(himin_i,12)) & -- 3
    CC(':') & -- 1
    CN(to_unsigned(himax_i,12)) & -- 3
    CC(' ') & -- 1
    CN(to_unsigned(vimin_i,12)) & -- 3
    CC(':') & -- 1
    CN(to_unsigned(vimax_i,12)) & -- 3
    CC(' ') & -- 1
    CN(to_unsigned(mire,4)) & -- 1
    CC(' ') & -- 1
    "1001" & iauto_n_i & -- 1
    "1001" & oauto_n_i & -- 1
    "1001" & inter & -- 1
    CS("          ") -- 10 
    ;
    
  ovo_in1<=
    CC(' ') & -- 1
    CN(to_unsigned(hmin_i,12)) & -- 3
    CC(':') & -- 1
    CN(to_unsigned(hmax_i,12)) & -- 3
    CC(' ') & -- 1
    CN(to_unsigned(vmin_i,12)) & -- 3
    CC(':') & -- 1
    CN(to_unsigned(vmax_i,12)) & -- 3
    CC(' ') & -- 1
    CS("               ") -- 15
    ;
  
  ovo_ena<='1'; -- Overlay
  
  ----------------------------------------------------------
  -- ROM / RAM

  reset_na<=NOT reset OR pll_locked;
  
END struct;
